// Copyright (c) 2018  LulinChen, All Rights Reserved
// AUTHOR : 	LulinChen
// AUTHOR'S EMAIL : lulinchen@aliyun.com 
// Release history
// VERSION Date AUTHOR DESCRIPTION

module rect0_rom(
	input 				clk,
	input		[11:0]	addr,
	output reg	[19:0]	q    // x y w h 5bit*4
	);
	reg					[19:0]	rom [4095:0];
	always @(posedge clk) q <= rom[addr];
	initial begin
		rom[ 0    ] = { 5'd6,	5'd4,	5'd12,	5'd9};
		rom[ 1    ] = { 5'd6,	5'd4,	5'd12,	5'd7};
		rom[ 2    ] = { 5'd3,	5'd9,	5'd18,	5'd9};
		rom[ 3    ] = { 5'd8,	5'd18,	5'd9,	5'd6};
		rom[ 4    ] = { 5'd3,	5'd5,	5'd4,	5'd19};
		rom[ 5    ] = { 5'd6,	5'd5,	5'd12,	5'd16};
		rom[ 6    ] = { 5'd5,	5'd8,	5'd12,	5'd6};
		rom[ 7    ] = { 5'd11,	5'd14,	5'd4,	5'd10};
		rom[ 8    ] = { 5'd4,	5'd0,	5'd7,	5'd6};
		rom[ 9    ] = { 5'd6,	5'd6,	5'd12,	5'd6};
		rom[ 10   ] = { 5'd6,	5'd4,	5'd12,	5'd7};
		rom[ 11   ] = { 5'd1,	5'd8,	5'd19,	5'd12};
		rom[ 12   ] = { 5'd0,	5'd2,	5'd24,	5'd3};
		rom[ 13   ] = { 5'd9,	5'd9,	5'd6,	5'd15};
		rom[ 14   ] = { 5'd5,	5'd6,	5'd14,	5'd10};
		rom[ 15   ] = { 5'd5,	5'd0,	5'd14,	5'd9};
		rom[ 16   ] = { 5'd13,	5'd11,	5'd9,	5'd6};
		rom[ 17   ] = { 5'd7,	5'd5,	5'd6,	5'd10};
		rom[ 18   ] = { 5'd10,	5'd8,	5'd6,	5'd10};
		rom[ 19   ] = { 5'd2,	5'd5,	5'd4,	5'd9};
		rom[ 20   ] = { 5'd18,	5'd0,	5'd6,	5'd11};
		rom[ 21   ] = { 5'd0,	5'd6,	5'd24,	5'd13};
		rom[ 22   ] = { 5'd9,	5'd6,	5'd6,	5'd9};
		rom[ 23   ] = { 5'd7,	5'd18,	5'd10,	5'd6};
		rom[ 24   ] = { 5'd5,	5'd7,	5'd14,	5'd12};
		rom[ 25   ] = { 5'd0,	5'd3,	5'd24,	5'd3};
		rom[ 26   ] = { 5'd5,	5'd8,	5'd15,	5'd6};
		rom[ 27   ] = { 5'd9,	5'd6,	5'd5,	5'd14};
		rom[ 28   ] = { 5'd9,	5'd5,	5'd6,	5'd10};
		rom[ 29   ] = { 5'd6,	5'd6,	5'd3,	5'd12};
		rom[ 30   ] = { 5'd3,	5'd21,	5'd18,	5'd3};
		rom[ 31   ] = { 5'd5,	5'd6,	5'd13,	5'd6};
		rom[ 32   ] = { 5'd18,	5'd1,	5'd6,	5'd15};
		rom[ 33   ] = { 5'd1,	5'd1,	5'd6,	5'd15};
		rom[ 34   ] = { 5'd0,	5'd8,	5'd24,	5'd15};
		rom[ 35   ] = { 5'd5,	5'd6,	5'd14,	5'd12};
		rom[ 36   ] = { 5'd2,	5'd12,	5'd21,	5'd12};
		rom[ 37   ] = { 5'd8,	5'd1,	5'd4,	5'd10};
		rom[ 38   ] = { 5'd2,	5'd13,	5'd20,	5'd10};
		rom[ 39   ] = { 5'd0,	5'd1,	5'd6,	5'd13};
		rom[ 40   ] = { 5'd20,	5'd2,	5'd4,	5'd13};
		rom[ 41   ] = { 5'd0,	5'd5,	5'd22,	5'd19};
		rom[ 42   ] = { 5'd18,	5'd4,	5'd6,	5'd9};
		rom[ 43   ] = { 5'd0,	5'd3,	5'd6,	5'd11};
		rom[ 44   ] = { 5'd12,	5'd1,	5'd4,	5'd9};
		rom[ 45   ] = { 5'd0,	5'd6,	5'd19,	5'd3};
		rom[ 46   ] = { 5'd12,	5'd1,	5'd4,	5'd9};
		rom[ 47   ] = { 5'd8,	5'd1,	5'd4,	5'd9};
		rom[ 48   ] = { 5'd5,	5'd5,	5'd14,	5'd14};
		rom[ 49   ] = { 5'd1,	5'd10,	5'd18,	5'd2};
		rom[ 50   ] = { 5'd17,	5'd13,	5'd4,	5'd11};
		rom[ 51   ] = { 5'd0,	5'd4,	5'd6,	5'd9};
		rom[ 52   ] = { 5'd6,	5'd4,	5'd12,	5'd9};
		rom[ 53   ] = { 5'd6,	5'd5,	5'd12,	5'd6};
		rom[ 54   ] = { 5'd0,	5'd1,	5'd24,	5'd5};
		rom[ 55   ] = { 5'd4,	5'd10,	5'd18,	5'd6};
		rom[ 56   ] = { 5'd2,	5'd17,	5'd12,	5'd6};
		rom[ 57   ] = { 5'd19,	5'd3,	5'd4,	5'd13};
		rom[ 58   ] = { 5'd1,	5'd3,	5'd4,	5'd13};
		rom[ 59   ] = { 5'd0,	5'd1,	5'd24,	5'd23};
		rom[ 60   ] = { 5'd1,	5'd7,	5'd8,	5'd12};
		rom[ 61   ] = { 5'd14,	5'd7,	5'd3,	5'd14};
		rom[ 62   ] = { 5'd3,	5'd12,	5'd16,	5'd6};
		rom[ 63   ] = { 5'd6,	5'd6,	5'd12,	5'd6};
		rom[ 64   ] = { 5'd8,	5'd7,	5'd6,	5'd12};
		rom[ 65   ] = { 5'd15,	5'd15,	5'd9,	5'd6};
		rom[ 66   ] = { 5'd1,	5'd17,	5'd18,	5'd3};
		rom[ 67   ] = { 5'd4,	5'd4,	5'd16,	5'd12};
		rom[ 68   ] = { 5'd0,	5'd1,	5'd4,	5'd20};
		rom[ 69   ] = { 5'd3,	5'd0,	5'd18,	5'd2};
		rom[ 70   ] = { 5'd1,	5'd5,	5'd20,	5'd14};
		rom[ 71   ] = { 5'd5,	5'd8,	5'd14,	5'd12};
		rom[ 72   ] = { 5'd3,	5'd14,	5'd7,	5'd9};
		rom[ 73   ] = { 5'd14,	5'd15,	5'd9,	5'd6};
		rom[ 74   ] = { 5'd1,	5'd15,	5'd9,	5'd6};
		rom[ 75   ] = { 5'd11,	5'd6,	5'd8,	5'd10};
		rom[ 76   ] = { 5'd5,	5'd5,	5'd14,	5'd14};
		rom[ 77   ] = { 5'd6,	5'd0,	5'd12,	5'd5};
		rom[ 78   ] = { 5'd9,	5'd0,	5'd6,	5'd9};
		rom[ 79   ] = { 5'd9,	5'd6,	5'd6,	5'd9};
		rom[ 80   ] = { 5'd7,	5'd0,	5'd6,	5'd9};
		rom[ 81   ] = { 5'd10,	5'd6,	5'd6,	5'd9};
		rom[ 82   ] = { 5'd8,	5'd6,	5'd6,	5'd9};
		rom[ 83   ] = { 5'd3,	5'd8,	5'd18,	5'd4};
		rom[ 84   ] = { 5'd6,	5'd0,	5'd12,	5'd9};
		rom[ 85   ] = { 5'd0,	5'd0,	5'd24,	5'd6};
		rom[ 86   ] = { 5'd4,	5'd7,	5'd16,	5'd12};
		rom[ 87   ] = { 5'd11,	5'd6,	5'd6,	5'd6};
		rom[ 88   ] = { 5'd0,	5'd20,	5'd24,	5'd3};
		rom[ 89   ] = { 5'd11,	5'd6,	5'd4,	5'd9};
		rom[ 90   ] = { 5'd4,	5'd13,	5'd15,	5'd4};
		rom[ 91   ] = { 5'd11,	5'd6,	5'd4,	5'd9};
		rom[ 92   ] = { 5'd9,	5'd6,	5'd4,	5'd9};
		rom[ 93   ] = { 5'd9,	5'd12,	5'd6,	5'd12};
		rom[ 94   ] = { 5'd1,	5'd22,	5'd18,	5'd2};
		rom[ 95   ] = { 5'd10,	5'd7,	5'd4,	5'd10};
		rom[ 96   ] = { 5'd6,	5'd7,	5'd8,	5'd10};
		rom[ 97   ] = { 5'd7,	5'd6,	5'd10,	5'd6};
		rom[ 98   ] = { 5'd0,	5'd14,	5'd10,	5'd4};
		rom[ 99   ] = { 5'd6,	5'd18,	5'd18,	5'd2};
		rom[ 100  ] = { 5'd1,	5'd1,	5'd22,	5'd3};
		rom[ 101  ] = { 5'd6,	5'd16,	5'd18,	5'd3};
		rom[ 102  ] = { 5'd2,	5'd4,	5'd6,	5'd15};
		rom[ 103  ] = { 5'd20,	5'd4,	5'd4,	5'd10};
		rom[ 104  ] = { 5'd0,	5'd4,	5'd4,	5'd10};
		rom[ 105  ] = { 5'd2,	5'd16,	5'd20,	5'd6};
		rom[ 106  ] = { 5'd0,	5'd12,	5'd8,	5'd9};
		rom[ 107  ] = { 5'd12,	5'd0,	5'd6,	5'd9};
		rom[ 108  ] = { 5'd5,	5'd10,	5'd6,	5'd6};
		rom[ 109  ] = { 5'd11,	5'd8,	5'd12,	5'd6};
		rom[ 110  ] = { 5'd0,	5'd8,	5'd12,	5'd6};
		rom[ 111  ] = { 5'd12,	5'd0,	5'd6,	5'd9};
		rom[ 112  ] = { 5'd6,	5'd0,	5'd6,	5'd9};
		rom[ 113  ] = { 5'd8,	5'd14,	5'd9,	5'd6};
		rom[ 114  ] = { 5'd0,	5'd16,	5'd9,	5'd6};
		rom[ 115  ] = { 5'd10,	5'd8,	5'd6,	5'd10};
		rom[ 116  ] = { 5'd3,	5'd19,	5'd12,	5'd3};
		rom[ 117  ] = { 5'd2,	5'd10,	5'd20,	5'd2};
		rom[ 118  ] = { 5'd2,	5'd9,	5'd18,	5'd12};
		rom[ 119  ] = { 5'd3,	5'd0,	5'd18,	5'd24};
		rom[ 120  ] = { 5'd5,	5'd6,	5'd14,	5'd10};
		rom[ 121  ] = { 5'd9,	5'd5,	5'd10,	5'd12};
		rom[ 122  ] = { 5'd4,	5'd5,	5'd12,	5'd12};
		rom[ 123  ] = { 5'd4,	5'd14,	5'd18,	5'd3};
		rom[ 124  ] = { 5'd6,	5'd13,	5'd8,	5'd8};
		rom[ 125  ] = { 5'd3,	5'd16,	5'd18,	5'd6};
		rom[ 126  ] = { 5'd0,	5'd0,	5'd6,	5'd6};
		rom[ 127  ] = { 5'd6,	5'd6,	5'd12,	5'd18};
		rom[ 128  ] = { 5'd6,	5'd1,	5'd4,	5'd14};
		rom[ 129  ] = { 5'd3,	5'd2,	5'd19,	5'd2};
		rom[ 130  ] = { 5'd1,	5'd8,	5'd22,	5'd13};
		rom[ 131  ] = { 5'd8,	5'd9,	5'd11,	5'd4};
		rom[ 132  ] = { 5'd0,	5'd12,	5'd15,	5'd10};
		rom[ 133  ] = { 5'd12,	5'd16,	5'd12,	5'd6};
		rom[ 134  ] = { 5'd0,	5'd16,	5'd12,	5'd6};
		rom[ 135  ] = { 5'd19,	5'd1,	5'd5,	5'd12};
		rom[ 136  ] = { 5'd0,	5'd2,	5'd24,	5'd4};
		rom[ 137  ] = { 5'd6,	5'd8,	5'd12,	5'd4};
		rom[ 138  ] = { 5'd7,	5'd5,	5'd9,	5'd6};
		rom[ 139  ] = { 5'd9,	5'd17,	5'd6,	5'd6};
		rom[ 140  ] = { 5'd0,	5'd7,	5'd22,	5'd15};
		rom[ 141  ] = { 5'd4,	5'd1,	5'd17,	5'd9};
		rom[ 142  ] = { 5'd7,	5'd5,	5'd6,	5'd10};
		rom[ 143  ] = { 5'd18,	5'd1,	5'd6,	5'd8};
		rom[ 144  ] = { 5'd0,	5'd1,	5'd6,	5'd7};
		rom[ 145  ] = { 5'd18,	5'd0,	5'd6,	5'd22};
		rom[ 146  ] = { 5'd0,	5'd0,	5'd6,	5'd22};
		rom[ 147  ] = { 5'd16,	5'd7,	5'd8,	5'd16};
		rom[ 148  ] = { 5'd2,	5'd10,	5'd19,	5'd6};
		rom[ 149  ] = { 5'd9,	5'd9,	5'd6,	5'd12};
		rom[ 150  ] = { 5'd2,	5'd15,	5'd17,	5'd6};
		rom[ 151  ] = { 5'd14,	5'd7,	5'd3,	5'd14};
		rom[ 152  ] = { 5'd5,	5'd6,	5'd8,	5'd10};
		rom[ 153  ] = { 5'd15,	5'd8,	5'd9,	5'd11};
		rom[ 154  ] = { 5'd0,	5'd8,	5'd9,	5'd11};
		rom[ 155  ] = { 5'd8,	5'd6,	5'd10,	5'd18};
		rom[ 156  ] = { 5'd7,	5'd7,	5'd3,	5'd14};
		rom[ 157  ] = { 5'd0,	5'd14,	5'd24,	5'd8};
		rom[ 158  ] = { 5'd1,	5'd10,	5'd18,	5'd14};
		rom[ 159  ] = { 5'd14,	5'd12,	5'd6,	5'd6};
		rom[ 160  ] = { 5'd7,	5'd0,	5'd10,	5'd16};
		rom[ 161  ] = { 5'd10,	5'd0,	5'd9,	5'd6};
		rom[ 162  ] = { 5'd4,	5'd3,	5'd16,	5'd4};
		rom[ 163  ] = { 5'd10,	5'd0,	5'd9,	5'd6};
		rom[ 164  ] = { 5'd1,	5'd1,	5'd20,	5'd4};
		rom[ 165  ] = { 5'd10,	5'd0,	5'd9,	5'd6};
		rom[ 166  ] = { 5'd5,	5'd0,	5'd9,	5'd6};
		rom[ 167  ] = { 5'd8,	5'd18,	5'd10,	5'd6};
		rom[ 168  ] = { 5'd6,	5'd3,	5'd6,	5'd9};
		rom[ 169  ] = { 5'd7,	5'd3,	5'd12,	5'd6};
		rom[ 170  ] = { 5'd0,	5'd10,	5'd18,	5'd3};
		rom[ 171  ] = { 5'd1,	5'd10,	5'd22,	5'd3};
		rom[ 172  ] = { 5'd5,	5'd11,	5'd8,	5'd8};
		rom[ 173  ] = { 5'd12,	5'd11,	5'd6,	5'd6};
		rom[ 174  ] = { 5'd6,	5'd11,	5'd6,	5'd6};
		rom[ 175  ] = { 5'd7,	5'd10,	5'd11,	5'd6};
		rom[ 176  ] = { 5'd0,	5'd13,	5'd24,	5'd4};
		rom[ 177  ] = { 5'd2,	5'd4,	5'd22,	5'd12};
		rom[ 178  ] = { 5'd2,	5'd0,	5'd20,	5'd17};
		rom[ 179  ] = { 5'd14,	5'd0,	5'd2,	5'd24};
		rom[ 180  ] = { 5'd8,	5'd0,	5'd2,	5'd24};
		rom[ 181  ] = { 5'd14,	5'd1,	5'd2,	5'd22};
		rom[ 182  ] = { 5'd8,	5'd1,	5'd2,	5'd22};
		rom[ 183  ] = { 5'd17,	5'd6,	5'd3,	5'd18};
		rom[ 184  ] = { 5'd6,	5'd14,	5'd9,	5'd6};
		rom[ 185  ] = { 5'd13,	5'd14,	5'd9,	5'd4};
		rom[ 186  ] = { 5'd3,	5'd18,	5'd18,	5'd3};
		rom[ 187  ] = { 5'd9,	5'd4,	5'd8,	5'd18};
		rom[ 188  ] = { 5'd0,	5'd17,	5'd18,	5'd3};
		rom[ 189  ] = { 5'd0,	5'd2,	5'd12,	5'd4};
		rom[ 190  ] = { 5'd6,	5'd8,	5'd14,	5'd6};
		rom[ 191  ] = { 5'd7,	5'd5,	5'd6,	5'd6};
		rom[ 192  ] = { 5'd10,	5'd5,	5'd6,	5'd16};
		rom[ 193  ] = { 5'd1,	5'd4,	5'd9,	5'd16};
		rom[ 194  ] = { 5'd5,	5'd0,	5'd18,	5'd9};
		rom[ 195  ] = { 5'd9,	5'd15,	5'd5,	5'd8};
		rom[ 196  ] = { 5'd20,	5'd0,	5'd4,	5'd9};
		rom[ 197  ] = { 5'd2,	5'd0,	5'd18,	5'd3};
		rom[ 198  ] = { 5'd5,	5'd22,	5'd19,	5'd2};
		rom[ 199  ] = { 5'd0,	5'd0,	5'd4,	5'd9};
		rom[ 200  ] = { 5'd5,	5'd6,	5'd19,	5'd18};
		rom[ 201  ] = { 5'd0,	5'd1,	5'd6,	5'd9};
		rom[ 202  ] = { 5'd6,	5'd5,	5'd14,	5'd12};
		rom[ 203  ] = { 5'd0,	5'd1,	5'd20,	5'd2};
		rom[ 204  ] = { 5'd1,	5'd2,	5'd22,	5'd3};
		rom[ 205  ] = { 5'd2,	5'd8,	5'd7,	5'd9};
		rom[ 206  ] = { 5'd2,	5'd12,	5'd22,	5'd4};
		rom[ 207  ] = { 5'd0,	5'd12,	5'd22,	5'd4};
		rom[ 208  ] = { 5'd9,	5'd7,	5'd6,	5'd11};
		rom[ 209  ] = { 5'd7,	5'd1,	5'd9,	5'd6};
		rom[ 210  ] = { 5'd11,	5'd2,	5'd4,	5'd10};
		rom[ 211  ] = { 5'd6,	5'd4,	5'd12,	5'd12};
		rom[ 212  ] = { 5'd18,	5'd1,	5'd6,	5'd15};
		rom[ 213  ] = { 5'd3,	5'd15,	5'd18,	5'd3};
		rom[ 214  ] = { 5'd18,	5'd5,	5'd6,	5'd9};
		rom[ 215  ] = { 5'd1,	5'd5,	5'd16,	5'd6};
		rom[ 216  ] = { 5'd11,	5'd0,	5'd6,	5'd9};
		rom[ 217  ] = { 5'd0,	5'd4,	5'd24,	5'd14};
		rom[ 218  ] = { 5'd13,	5'd0,	5'd4,	5'd13};
		rom[ 219  ] = { 5'd7,	5'd0,	5'd4,	5'd13};
		rom[ 220  ] = { 5'd11,	5'd6,	5'd6,	5'd9};
		rom[ 221  ] = { 5'd8,	5'd7,	5'd6,	5'd9};
		rom[ 222  ] = { 5'd13,	5'd17,	5'd9,	5'd6};
		rom[ 223  ] = { 5'd2,	5'd18,	5'd14,	5'd6};
		rom[ 224  ] = { 5'd3,	5'd18,	5'd18,	5'd4};
		rom[ 225  ] = { 5'd0,	5'd20,	5'd15,	5'd4};
		rom[ 226  ] = { 5'd9,	5'd15,	5'd15,	5'd9};
		rom[ 227  ] = { 5'd4,	5'd4,	5'd16,	5'd4};
		rom[ 228  ] = { 5'd7,	5'd6,	5'd10,	5'd6};
		rom[ 229  ] = { 5'd0,	5'd14,	5'd15,	5'd10};
		rom[ 230  ] = { 5'd7,	5'd9,	5'd10,	5'd14};
		rom[ 231  ] = { 5'd7,	5'd6,	5'd6,	5'd9};
		rom[ 232  ] = { 5'd3,	5'd6,	5'd18,	5'd3};
		rom[ 233  ] = { 5'd0,	5'd10,	5'd18,	5'd3};
		rom[ 234  ] = { 5'd3,	5'd16,	5'd18,	5'd4};
		rom[ 235  ] = { 5'd4,	5'd6,	5'd14,	5'd6};
		rom[ 236  ] = { 5'd13,	5'd0,	5'd2,	5'd18};
		rom[ 237  ] = { 5'd9,	5'd0,	5'd2,	5'd18};
		rom[ 238  ] = { 5'd5,	5'd7,	5'd15,	5'd10};
		rom[ 239  ] = { 5'd1,	5'd20,	5'd21,	5'd4};
		rom[ 240  ] = { 5'd10,	5'd5,	5'd5,	5'd18};
		rom[ 241  ] = { 5'd0,	5'd2,	5'd24,	5'd6};
		rom[ 242  ] = { 5'd1,	5'd1,	5'd22,	5'd8};
		rom[ 243  ] = { 5'd4,	5'd0,	5'd15,	5'd9};
		rom[ 244  ] = { 5'd0,	5'd0,	5'd24,	5'd19};
		rom[ 245  ] = { 5'd2,	5'd21,	5'd18,	5'd3};
		rom[ 246  ] = { 5'd9,	5'd7,	5'd10,	5'd4};
		rom[ 247  ] = { 5'd5,	5'd7,	5'd10,	5'd4};
		rom[ 248  ] = { 5'd17,	5'd8,	5'd6,	5'd16};
		rom[ 249  ] = { 5'd1,	5'd15,	5'd20,	5'd4};
		rom[ 250  ] = { 5'd14,	5'd15,	5'd10,	5'd6};
		rom[ 251  ] = { 5'd3,	5'd0,	5'd16,	5'd9};
		rom[ 252  ] = { 5'd15,	5'd6,	5'd7,	5'd15};
		rom[ 253  ] = { 5'd9,	5'd1,	5'd6,	5'd13};
		rom[ 254  ] = { 5'd17,	5'd2,	5'd6,	5'd14};
		rom[ 255  ] = { 5'd3,	5'd14,	5'd12,	5'd10};
		rom[ 256  ] = { 5'd7,	5'd6,	5'd10,	5'd6};
		rom[ 257  ] = { 5'd1,	5'd2,	5'd6,	5'd14};
		rom[ 258  ] = { 5'd10,	5'd4,	5'd5,	5'd12};
		rom[ 259  ] = { 5'd0,	5'd17,	5'd24,	5'd5};
		rom[ 260  ] = { 5'd15,	5'd7,	5'd5,	5'd12};
		rom[ 261  ] = { 5'd3,	5'd1,	5'd6,	5'd12};
		rom[ 262  ] = { 5'd12,	5'd13,	5'd6,	5'd6};
		rom[ 263  ] = { 5'd6,	5'd13,	5'd6,	5'd6};
		rom[ 264  ] = { 5'd14,	5'd6,	5'd3,	5'd16};
		rom[ 265  ] = { 5'd1,	5'd12,	5'd13,	5'd6};
		rom[ 266  ] = { 5'd13,	5'd1,	5'd4,	5'd9};
		rom[ 267  ] = { 5'd7,	5'd0,	5'd9,	5'd6};
		rom[ 268  ] = { 5'd12,	5'd2,	5'd6,	5'd9};
		rom[ 269  ] = { 5'd6,	5'd2,	5'd6,	5'd9};
		rom[ 270  ] = { 5'd6,	5'd18,	5'd12,	5'd6};
		rom[ 271  ] = { 5'd7,	5'd6,	5'd6,	5'd9};
		rom[ 272  ] = { 5'd7,	5'd7,	5'd12,	5'd3};
		rom[ 273  ] = { 5'd8,	5'd3,	5'd8,	5'd21};
		rom[ 274  ] = { 5'd7,	5'd4,	5'd10,	5'd12};
		rom[ 275  ] = { 5'd0,	5'd1,	5'd6,	5'd9};
		rom[ 276  ] = { 5'd15,	5'd2,	5'd2,	5'd20};
		rom[ 277  ] = { 5'd0,	5'd3,	5'd6,	5'd9};
		rom[ 278  ] = { 5'd15,	5'd3,	5'd2,	5'd21};
		rom[ 279  ] = { 5'd7,	5'd0,	5'd2,	5'd23};
		rom[ 280  ] = { 5'd15,	5'd8,	5'd9,	5'd4};
		rom[ 281  ] = { 5'd0,	5'd8,	5'd9,	5'd4};
		rom[ 282  ] = { 5'd8,	5'd14,	5'd9,	5'd6};
		rom[ 283  ] = { 5'd0,	5'd14,	5'd9,	5'd6};
		rom[ 284  ] = { 5'd3,	5'd10,	5'd18,	5'd4};
		rom[ 285  ] = { 5'd0,	5'd0,	5'd24,	5'd19};
		rom[ 286  ] = { 5'd9,	5'd1,	5'd8,	5'd12};
		rom[ 287  ] = { 5'd10,	5'd6,	5'd4,	5'd10};
		rom[ 288  ] = { 5'd7,	5'd9,	5'd10,	5'd12};
		rom[ 289  ] = { 5'd5,	5'd0,	5'd3,	5'd19};
		rom[ 290  ] = { 5'd14,	5'd0,	5'd6,	5'd10};
		rom[ 291  ] = { 5'd2,	5'd0,	5'd6,	5'd12};
		rom[ 292  ] = { 5'd0,	5'd11,	5'd24,	5'd2};
		rom[ 293  ] = { 5'd4,	5'd9,	5'd13,	5'd4};
		rom[ 294  ] = { 5'd9,	5'd8,	5'd6,	5'd9};
		rom[ 295  ] = { 5'd0,	5'd12,	5'd16,	5'd4};
		rom[ 296  ] = { 5'd18,	5'd12,	5'd6,	5'd9};
		rom[ 297  ] = { 5'd0,	5'd12,	5'd6,	5'd9};
		rom[ 298  ] = { 5'd8,	5'd7,	5'd10,	5'd4};
		rom[ 299  ] = { 5'd8,	5'd7,	5'd6,	5'd9};
		rom[ 300  ] = { 5'd11,	5'd0,	5'd6,	5'd9};
		rom[ 301  ] = { 5'd7,	5'd0,	5'd6,	5'd9};
		rom[ 302  ] = { 5'd12,	5'd3,	5'd6,	5'd15};
		rom[ 303  ] = { 5'd6,	5'd3,	5'd6,	5'd15};
		rom[ 304  ] = { 5'd15,	5'd2,	5'd9,	5'd4};
		rom[ 305  ] = { 5'd5,	5'd10,	5'd6,	5'd7};
		rom[ 306  ] = { 5'd9,	5'd14,	5'd6,	5'd10};
		rom[ 307  ] = { 5'd7,	5'd13,	5'd5,	5'd8};
		rom[ 308  ] = { 5'd14,	5'd5,	5'd3,	5'd16};
		rom[ 309  ] = { 5'd2,	5'd17,	5'd18,	5'd3};
		rom[ 310  ] = { 5'd5,	5'd18,	5'd19,	5'd3};
		rom[ 311  ] = { 5'd9,	5'd0,	5'd6,	5'd9};
		rom[ 312  ] = { 5'd12,	5'd4,	5'd3,	5'd18};
		rom[ 313  ] = { 5'd9,	5'd4,	5'd3,	5'd18};
		rom[ 314  ] = { 5'd3,	5'd3,	5'd18,	5'd9};
		rom[ 315  ] = { 5'd6,	5'd1,	5'd6,	5'd14};
		rom[ 316  ] = { 5'd12,	5'd16,	5'd9,	5'd6};
		rom[ 317  ] = { 5'd1,	5'd3,	5'd20,	5'd16};
		rom[ 318  ] = { 5'd12,	5'd5,	5'd6,	5'd12};
		rom[ 319  ] = { 5'd1,	5'd2,	5'd22,	5'd16};
		rom[ 320  ] = { 5'd10,	5'd14,	5'd5,	5'd10};
		rom[ 321  ] = { 5'd3,	5'd21,	5'd18,	5'd3};
		rom[ 322  ] = { 5'd10,	5'd14,	5'd6,	5'd10};
		rom[ 323  ] = { 5'd0,	5'd2,	5'd24,	5'd4};
		rom[ 324  ] = { 5'd6,	5'd4,	5'd12,	5'd9};
		rom[ 325  ] = { 5'd6,	5'd6,	5'd12,	5'd5};
		rom[ 326  ] = { 5'd5,	5'd8,	5'd14,	5'd12};
		rom[ 327  ] = { 5'd4,	5'd14,	5'd8,	5'd10};
		rom[ 328  ] = { 5'd11,	5'd6,	5'd5,	5'd14};
		rom[ 329  ] = { 5'd7,	5'd6,	5'd3,	5'd16};
		rom[ 330  ] = { 5'd3,	5'd7,	5'd18,	5'd8};
		rom[ 331  ] = { 5'd2,	5'd3,	5'd20,	5'd2};
		rom[ 332  ] = { 5'd3,	5'd12,	5'd19,	5'd6};
		rom[ 333  ] = { 5'd8,	5'd6,	5'd6,	5'd9};
		rom[ 334  ] = { 5'd16,	5'd6,	5'd6,	5'd14};
		rom[ 335  ] = { 5'd7,	5'd9,	5'd6,	5'd12};
		rom[ 336  ] = { 5'd18,	5'd6,	5'd6,	5'd18};
		rom[ 337  ] = { 5'd0,	5'd6,	5'd6,	5'd18};
		rom[ 338  ] = { 5'd18,	5'd2,	5'd6,	5'd9};
		rom[ 339  ] = { 5'd3,	5'd18,	5'd15,	5'd6};
		rom[ 340  ] = { 5'd18,	5'd2,	5'd6,	5'd9};
		rom[ 341  ] = { 5'd0,	5'd2,	5'd6,	5'd9};
		rom[ 342  ] = { 5'd5,	5'd10,	5'd18,	5'd2};
		rom[ 343  ] = { 5'd6,	5'd0,	5'd12,	5'd6};
		rom[ 344  ] = { 5'd10,	5'd0,	5'd6,	5'd9};
		rom[ 345  ] = { 5'd8,	5'd0,	5'd6,	5'd9};
		rom[ 346  ] = { 5'd15,	5'd12,	5'd9,	5'd6};
		rom[ 347  ] = { 5'd3,	5'd6,	5'd13,	5'd6};
		rom[ 348  ] = { 5'd15,	5'd12,	5'd9,	5'd6};
		rom[ 349  ] = { 5'd2,	5'd5,	5'd6,	5'd15};
		rom[ 350  ] = { 5'd8,	5'd8,	5'd9,	5'd6};
		rom[ 351  ] = { 5'd8,	5'd6,	5'd3,	5'd14};
		rom[ 352  ] = { 5'd15,	5'd12,	5'd9,	5'd6};
		rom[ 353  ] = { 5'd4,	5'd12,	5'd10,	5'd4};
		rom[ 354  ] = { 5'd13,	5'd1,	5'd4,	5'd19};
		rom[ 355  ] = { 5'd7,	5'd1,	5'd4,	5'd19};
		rom[ 356  ] = { 5'd18,	5'd9,	5'd6,	5'd9};
		rom[ 357  ] = { 5'd1,	5'd21,	5'd18,	5'd3};
		rom[ 358  ] = { 5'd14,	5'd13,	5'd10,	5'd9};
		rom[ 359  ] = { 5'd1,	5'd13,	5'd22,	5'd4};
		rom[ 360  ] = { 5'd4,	5'd6,	5'd16,	5'd6};
		rom[ 361  ] = { 5'd1,	5'd0,	5'd18,	5'd22};
		rom[ 362  ] = { 5'd10,	5'd7,	5'd8,	5'd14};
		rom[ 363  ] = { 5'd0,	5'd4,	5'd6,	5'd20};
		rom[ 364  ] = { 5'd15,	5'd0,	5'd6,	5'd9};
		rom[ 365  ] = { 5'd3,	5'd0,	5'd6,	5'd9};
		rom[ 366  ] = { 5'd15,	5'd12,	5'd6,	5'd12};
		rom[ 367  ] = { 5'd3,	5'd12,	5'd6,	5'd12};
		rom[ 368  ] = { 5'd15,	5'd12,	5'd9,	5'd6};
		rom[ 369  ] = { 5'd0,	5'd12,	5'd9,	5'd6};
		rom[ 370  ] = { 5'd4,	5'd14,	5'd19,	5'd3};
		rom[ 371  ] = { 5'd2,	5'd13,	5'd19,	5'd3};
		rom[ 372  ] = { 5'd14,	5'd15,	5'd10,	5'd6};
		rom[ 373  ] = { 5'd6,	5'd0,	5'd10,	5'd12};
		rom[ 374  ] = { 5'd17,	5'd1,	5'd6,	5'd12};
		rom[ 375  ] = { 5'd1,	5'd1,	5'd6,	5'd12};
		rom[ 376  ] = { 5'd16,	5'd14,	5'd6,	5'd9};
		rom[ 377  ] = { 5'd7,	5'd3,	5'd9,	5'd12};
		rom[ 378  ] = { 5'd12,	5'd1,	5'd4,	5'd12};
		rom[ 379  ] = { 5'd4,	5'd0,	5'd14,	5'd8};
		rom[ 380  ] = { 5'd10,	5'd6,	5'd6,	5'd9};
		rom[ 381  ] = { 5'd2,	5'd10,	5'd18,	5'd3};
		rom[ 382  ] = { 5'd15,	5'd15,	5'd9,	5'd6};
		rom[ 383  ] = { 5'd0,	5'd1,	5'd21,	5'd23};
		rom[ 384  ] = { 5'd6,	5'd9,	5'd17,	5'd4};
		rom[ 385  ] = { 5'd1,	5'd0,	5'd11,	5'd18};
		rom[ 386  ] = { 5'd6,	5'd15,	5'd13,	5'd6};
		rom[ 387  ] = { 5'd0,	5'd15,	5'd9,	5'd6};
		rom[ 388  ] = { 5'd8,	5'd7,	5'd15,	5'd4};
		rom[ 389  ] = { 5'd9,	5'd12,	5'd6,	5'd9};
		rom[ 390  ] = { 5'd6,	5'd8,	5'd18,	5'd3};
		rom[ 391  ] = { 5'd0,	5'd14,	5'd24,	5'd4};
		rom[ 392  ] = { 5'd16,	5'd10,	5'd3,	5'd12};
		rom[ 393  ] = { 5'd0,	5'd3,	5'd24,	5'd3};
		rom[ 394  ] = { 5'd14,	5'd17,	5'd10,	5'd6};
		rom[ 395  ] = { 5'd1,	5'd13,	5'd18,	5'd3};
		rom[ 396  ] = { 5'd5,	5'd0,	5'd18,	5'd9};
		rom[ 397  ] = { 5'd4,	5'd3,	5'd16,	5'd9};
		rom[ 398  ] = { 5'd16,	5'd5,	5'd3,	5'd12};
		rom[ 399  ] = { 5'd0,	5'd7,	5'd18,	5'd4};
		rom[ 400  ] = { 5'd10,	5'd6,	5'd6,	5'd9};
		rom[ 401  ] = { 5'd9,	5'd8,	5'd6,	5'd10};
		rom[ 402  ] = { 5'd9,	5'd15,	5'd6,	5'd9};
		rom[ 403  ] = { 5'd3,	5'd1,	5'd18,	5'd21};
		rom[ 404  ] = { 5'd6,	5'd8,	5'd12,	5'd7};
		rom[ 405  ] = { 5'd8,	5'd5,	5'd6,	5'd9};
		rom[ 406  ] = { 5'd0,	5'd2,	5'd24,	5'd4};
		rom[ 407  ] = { 5'd14,	5'd7,	5'd5,	5'd12};
		rom[ 408  ] = { 5'd5,	5'd7,	5'd5,	5'd12};
		rom[ 409  ] = { 5'd9,	5'd6,	5'd6,	5'd9};
		rom[ 410  ] = { 5'd0,	5'd1,	5'd6,	5'd17};
		rom[ 411  ] = { 5'd3,	5'd1,	5'd19,	5'd9};
		rom[ 412  ] = { 5'd3,	5'd18,	5'd12,	5'd6};
		rom[ 413  ] = { 5'd20,	5'd4,	5'd4,	5'd19};
		rom[ 414  ] = { 5'd0,	5'd16,	5'd10,	5'd7};
		rom[ 415  ] = { 5'd8,	5'd7,	5'd10,	5'd12};
		rom[ 416  ] = { 5'd6,	5'd7,	5'd10,	5'd12};
		rom[ 417  ] = { 5'd9,	5'd2,	5'd9,	5'd6};
		rom[ 418  ] = { 5'd1,	5'd20,	5'd21,	5'd4};
		rom[ 419  ] = { 5'd9,	5'd12,	5'd9,	5'd6};
		rom[ 420  ] = { 5'd7,	5'd2,	5'd9,	5'd6};
		rom[ 421  ] = { 5'd13,	5'd0,	5'd4,	5'd14};
		rom[ 422  ] = { 5'd7,	5'd0,	5'd4,	5'd14};
		rom[ 423  ] = { 5'd14,	5'd15,	5'd9,	5'd6};
		rom[ 424  ] = { 5'd2,	5'd8,	5'd18,	5'd5};
		rom[ 425  ] = { 5'd18,	5'd3,	5'd6,	5'd11};
		rom[ 426  ] = { 5'd6,	5'd5,	5'd11,	5'd14};
		rom[ 427  ] = { 5'd18,	5'd4,	5'd6,	5'd9};
		rom[ 428  ] = { 5'd7,	5'd6,	5'd9,	5'd6};
		rom[ 429  ] = { 5'd18,	5'd4,	5'd6,	5'd9};
		rom[ 430  ] = { 5'd0,	5'd4,	5'd6,	5'd9};
		rom[ 431  ] = { 5'd9,	5'd4,	5'd9,	5'd4};
		rom[ 432  ] = { 5'd0,	5'd22,	5'd19,	5'd2};
		rom[ 433  ] = { 5'd17,	5'd14,	5'd6,	5'd9};
		rom[ 434  ] = { 5'd1,	5'd14,	5'd6,	5'd9};
		rom[ 435  ] = { 5'd14,	5'd11,	5'd4,	5'd9};
		rom[ 436  ] = { 5'd6,	5'd11,	5'd4,	5'd9};
		rom[ 437  ] = { 5'd3,	5'd9,	5'd18,	5'd7};
		rom[ 438  ] = { 5'd9,	5'd12,	5'd6,	5'd10};
		rom[ 439  ] = { 5'd12,	5'd0,	5'd6,	5'd9};
		rom[ 440  ] = { 5'd6,	5'd0,	5'd6,	5'd9};
		rom[ 441  ] = { 5'd6,	5'd17,	5'd18,	5'd3};
		rom[ 442  ] = { 5'd1,	5'd17,	5'd18,	5'd3};
		rom[ 443  ] = { 5'd10,	5'd6,	5'd11,	5'd12};
		rom[ 444  ] = { 5'd5,	5'd6,	5'd14,	5'd6};
		rom[ 445  ] = { 5'd5,	5'd4,	5'd15,	5'd4};
		rom[ 446  ] = { 5'd0,	5'd0,	5'd22,	5'd2};
		rom[ 447  ] = { 5'd0,	5'd0,	5'd24,	5'd24};
		rom[ 448  ] = { 5'd1,	5'd15,	5'd18,	5'd4};
		rom[ 449  ] = { 5'd6,	5'd8,	5'd12,	5'd9};
		rom[ 450  ] = { 5'd4,	5'd12,	5'd7,	5'd12};
		rom[ 451  ] = { 5'd1,	5'd2,	5'd22,	5'd6};
		rom[ 452  ] = { 5'd5,	5'd20,	5'd14,	5'd3};
		rom[ 453  ] = { 5'd0,	5'd0,	5'd24,	5'd16};
		rom[ 454  ] = { 5'd3,	5'd13,	5'd18,	5'd4};
		rom[ 455  ] = { 5'd2,	5'd10,	5'd22,	5'd2};
		rom[ 456  ] = { 5'd6,	5'd3,	5'd11,	5'd8};
		rom[ 457  ] = { 5'd14,	5'd5,	5'd6,	5'd6};
		rom[ 458  ] = { 5'd0,	5'd7,	5'd24,	5'd6};
		rom[ 459  ] = { 5'd14,	5'd0,	5'd10,	5'd10};
		rom[ 460  ] = { 5'd0,	5'd0,	5'd10,	5'd10};
		rom[ 461  ] = { 5'd0,	5'd1,	5'd24,	5'd4};
		rom[ 462  ] = { 5'd0,	5'd17,	5'd18,	5'd3};
		rom[ 463  ] = { 5'd5,	5'd15,	5'd16,	5'd6};
		rom[ 464  ] = { 5'd3,	5'd15,	5'd16,	5'd6};
		rom[ 465  ] = { 5'd6,	5'd16,	5'd18,	5'd3};
		rom[ 466  ] = { 5'd0,	5'd13,	5'd21,	5'd10};
		rom[ 467  ] = { 5'd13,	5'd0,	5'd6,	5'd24};
		rom[ 468  ] = { 5'd7,	5'd4,	5'd6,	5'd11};
		rom[ 469  ] = { 5'd9,	5'd5,	5'd9,	5'd6};
		rom[ 470  ] = { 5'd1,	5'd4,	5'd2,	5'd20};
		rom[ 471  ] = { 5'd13,	5'd0,	5'd6,	5'd24};
		rom[ 472  ] = { 5'd5,	5'd0,	5'd6,	5'd24};
		rom[ 473  ] = { 5'd16,	5'd7,	5'd6,	5'd14};
		rom[ 474  ] = { 5'd4,	5'd7,	5'd4,	5'd12};
		rom[ 475  ] = { 5'd0,	5'd5,	5'd24,	5'd14};
		rom[ 476  ] = { 5'd5,	5'd13,	5'd10,	5'd6};
		rom[ 477  ] = { 5'd12,	5'd0,	5'd6,	5'd9};
		rom[ 478  ] = { 5'd2,	5'd7,	5'd6,	5'd14};
		rom[ 479  ] = { 5'd15,	5'd2,	5'd9,	5'd15};
		rom[ 480  ] = { 5'd0,	5'd2,	5'd6,	5'd9};
		rom[ 481  ] = { 5'd12,	5'd2,	5'd10,	5'd14};
		rom[ 482  ] = { 5'd11,	5'd6,	5'd2,	5'd18};
		rom[ 483  ] = { 5'd9,	5'd5,	5'd15,	5'd6};
		rom[ 484  ] = { 5'd8,	5'd6,	5'd6,	5'd10};
		rom[ 485  ] = { 5'd12,	5'd0,	5'd6,	5'd9};
		rom[ 486  ] = { 5'd3,	5'd3,	5'd9,	5'd7};
		rom[ 487  ] = { 5'd6,	5'd7,	5'd14,	5'd3};
		rom[ 488  ] = { 5'd7,	5'd7,	5'd8,	5'd6};
		rom[ 489  ] = { 5'd12,	5'd7,	5'd7,	5'd12};
		rom[ 490  ] = { 5'd10,	5'd6,	5'd4,	5'd18};
		rom[ 491  ] = { 5'd16,	5'd14,	5'd6,	5'd9};
		rom[ 492  ] = { 5'd4,	5'd0,	5'd6,	5'd13};
		rom[ 493  ] = { 5'd2,	5'd2,	5'd21,	5'd3};
		rom[ 494  ] = { 5'd5,	5'd4,	5'd5,	5'd12};
		rom[ 495  ] = { 5'd10,	5'd3,	5'd4,	5'd10};
		rom[ 496  ] = { 5'd8,	5'd4,	5'd5,	5'd8};
		rom[ 497  ] = { 5'd6,	5'd0,	5'd11,	5'd9};
		rom[ 498  ] = { 5'd6,	5'd6,	5'd12,	5'd5};
		rom[ 499  ] = { 5'd0,	5'd0,	5'd24,	5'd5};
		rom[ 500  ] = { 5'd1,	5'd10,	5'd23,	5'd6};
		rom[ 501  ] = { 5'd3,	5'd21,	5'd18,	5'd3};
		rom[ 502  ] = { 5'd3,	5'd6,	5'd21,	5'd6};
		rom[ 503  ] = { 5'd0,	5'd5,	5'd6,	5'd12};
		rom[ 504  ] = { 5'd10,	5'd2,	5'd4,	5'd15};
		rom[ 505  ] = { 5'd8,	5'd7,	5'd8,	5'd10};
		rom[ 506  ] = { 5'd5,	5'd7,	5'd15,	5'd12};
		rom[ 507  ] = { 5'd0,	5'd17,	5'd10,	5'd6};
		rom[ 508  ] = { 5'd14,	5'd18,	5'd9,	5'd6};
		rom[ 509  ] = { 5'd9,	5'd6,	5'd6,	5'd16};
		rom[ 510  ] = { 5'd14,	5'd18,	5'd9,	5'd6};
		rom[ 511  ] = { 5'd1,	5'd18,	5'd9,	5'd6};
		rom[ 512  ] = { 5'd15,	5'd9,	5'd9,	5'd6};
		rom[ 513  ] = { 5'd0,	5'd9,	5'd9,	5'd6};
		rom[ 514  ] = { 5'd17,	5'd3,	5'd6,	5'd9};
		rom[ 515  ] = { 5'd2,	5'd17,	5'd18,	5'd3};
		rom[ 516  ] = { 5'd3,	5'd15,	5'd21,	5'd6};
		rom[ 517  ] = { 5'd9,	5'd17,	5'd6,	5'd6};
		rom[ 518  ] = { 5'd18,	5'd3,	5'd6,	5'd9};
		rom[ 519  ] = { 5'd0,	5'd3,	5'd6,	5'd9};
		rom[ 520  ] = { 5'd4,	5'd0,	5'd16,	5'd10};
		rom[ 521  ] = { 5'd2,	5'd0,	5'd10,	5'd16};
		rom[ 522  ] = { 5'd14,	5'd0,	5'd10,	5'd5};
		rom[ 523  ] = { 5'd0,	5'd0,	5'd10,	5'd5};
		rom[ 524  ] = { 5'd18,	5'd3,	5'd6,	5'd10};
		rom[ 525  ] = { 5'd5,	5'd11,	5'd12,	5'd6};
		rom[ 526  ] = { 5'd21,	5'd0,	5'd3,	5'd18};
		rom[ 527  ] = { 5'd6,	5'd0,	5'd6,	5'd9};
		rom[ 528  ] = { 5'd8,	5'd8,	5'd9,	5'd7};
		rom[ 529  ] = { 5'd7,	5'd12,	5'd8,	5'd10};
		rom[ 530  ] = { 5'd21,	5'd0,	5'd3,	5'd18};
		rom[ 531  ] = { 5'd10,	5'd6,	5'd4,	5'd9};
		rom[ 532  ] = { 5'd15,	5'd0,	5'd9,	5'd6};
		rom[ 533  ] = { 5'd0,	5'd2,	5'd24,	5'd3};
		rom[ 534  ] = { 5'd11,	5'd7,	5'd6,	5'd9};
		rom[ 535  ] = { 5'd7,	5'd6,	5'd6,	5'd10};
		rom[ 536  ] = { 5'd12,	5'd1,	5'd6,	5'd12};
		rom[ 537  ] = { 5'd6,	5'd4,	5'd12,	5'd12};
		rom[ 538  ] = { 5'd14,	5'd3,	5'd2,	5'd21};
		rom[ 539  ] = { 5'd6,	5'd1,	5'd12,	5'd8};
		rom[ 540  ] = { 5'd3,	5'd0,	5'd18,	5'd8};
		rom[ 541  ] = { 5'd3,	5'd0,	5'd18,	5'd3};
		rom[ 542  ] = { 5'd0,	5'd13,	5'd24,	5'd4};
		rom[ 543  ] = { 5'd10,	5'd5,	5'd4,	5'd9};
		rom[ 544  ] = { 5'd11,	5'd1,	5'd6,	5'd9};
		rom[ 545  ] = { 5'd6,	5'd2,	5'd6,	5'd22};
		rom[ 546  ] = { 5'd16,	5'd10,	5'd8,	5'd14};
		rom[ 547  ] = { 5'd3,	5'd4,	5'd16,	5'd15};
		rom[ 548  ] = { 5'd16,	5'd10,	5'd8,	5'd14};
		rom[ 549  ] = { 5'd0,	5'd10,	5'd8,	5'd14};
		rom[ 550  ] = { 5'd10,	5'd14,	5'd11,	5'd6};
		rom[ 551  ] = { 5'd0,	5'd7,	5'd24,	5'd9};
		rom[ 552  ] = { 5'd13,	5'd1,	5'd4,	5'd16};
		rom[ 553  ] = { 5'd7,	5'd1,	5'd4,	5'd16};
		rom[ 554  ] = { 5'd5,	5'd5,	5'd16,	5'd8};
		rom[ 555  ] = { 5'd0,	5'd9,	5'd6,	5'd9};
		rom[ 556  ] = { 5'd6,	5'd16,	5'd18,	5'd3};
		rom[ 557  ] = { 5'd3,	5'd12,	5'd6,	5'd9};
		rom[ 558  ] = { 5'd8,	5'd14,	5'd9,	5'd6};
		rom[ 559  ] = { 5'd2,	5'd13,	5'd8,	5'd10};
		rom[ 560  ] = { 5'd15,	5'd5,	5'd3,	5'd18};
		rom[ 561  ] = { 5'd3,	5'd5,	5'd18,	5'd3};
		rom[ 562  ] = { 5'd17,	5'd5,	5'd6,	5'd11};
		rom[ 563  ] = { 5'd1,	5'd5,	5'd6,	5'd11};
		rom[ 564  ] = { 5'd19,	5'd1,	5'd4,	5'd9};
		rom[ 565  ] = { 5'd1,	5'd1,	5'd4,	5'd9};
		rom[ 566  ] = { 5'd4,	5'd15,	5'd18,	5'd9};
		rom[ 567  ] = { 5'd6,	5'd9,	5'd12,	5'd4};
		rom[ 568  ] = { 5'd15,	5'd2,	5'd9,	5'd6};
		rom[ 569  ] = { 5'd0,	5'd2,	5'd9,	5'd6};
		rom[ 570  ] = { 5'd15,	5'd0,	5'd6,	5'd17};
		rom[ 571  ] = { 5'd3,	5'd0,	5'd6,	5'd17};
		rom[ 572  ] = { 5'd8,	5'd17,	5'd9,	5'd4};
		rom[ 573  ] = { 5'd6,	5'd5,	5'd3,	5'd18};
		rom[ 574  ] = { 5'd5,	5'd2,	5'd14,	5'd12};
		rom[ 575  ] = { 5'd10,	5'd2,	5'd3,	5'd12};
		rom[ 576  ] = { 5'd10,	5'd7,	5'd14,	5'd15};
		rom[ 577  ] = { 5'd0,	5'd7,	5'd14,	5'd15};
		rom[ 578  ] = { 5'd15,	5'd0,	5'd9,	5'd6};
		rom[ 579  ] = { 5'd0,	5'd0,	5'd9,	5'd6};
		rom[ 580  ] = { 5'd12,	5'd6,	5'd6,	5'd14};
		rom[ 581  ] = { 5'd9,	5'd7,	5'd6,	5'd9};
		rom[ 582  ] = { 5'd12,	5'd6,	5'd6,	5'd15};
		rom[ 583  ] = { 5'd6,	5'd6,	5'd6,	5'd15};
		rom[ 584  ] = { 5'd15,	5'd3,	5'd8,	5'd9};
		rom[ 585  ] = { 5'd0,	5'd0,	5'd9,	5'd21};
		rom[ 586  ] = { 5'd11,	5'd9,	5'd8,	5'd12};
		rom[ 587  ] = { 5'd6,	5'd7,	5'd10,	5'd12};
		rom[ 588  ] = { 5'd10,	5'd6,	5'd4,	5'd18};
		rom[ 589  ] = { 5'd0,	5'd0,	5'd6,	5'd9};
		rom[ 590  ] = { 5'd3,	5'd14,	5'd18,	5'd3};
		rom[ 591  ] = { 5'd3,	5'd14,	5'd8,	5'd10};
		rom[ 592  ] = { 5'd0,	5'd12,	5'd24,	5'd4};
		rom[ 593  ] = { 5'd0,	5'd2,	5'd3,	5'd20};
		rom[ 594  ] = { 5'd12,	5'd16,	5'd10,	5'd8};
		rom[ 595  ] = { 5'd2,	5'd16,	5'd10,	5'd8};
		rom[ 596  ] = { 5'd7,	5'd0,	5'd10,	5'd9};
		rom[ 597  ] = { 5'd0,	5'd0,	5'd24,	5'd3};
		rom[ 598  ] = { 5'd3,	5'd8,	5'd15,	5'd4};
		rom[ 599  ] = { 5'd6,	5'd5,	5'd12,	5'd6};
		rom[ 600  ] = { 5'd5,	5'd13,	5'd14,	5'd6};
		rom[ 601  ] = { 5'd11,	5'd14,	5'd4,	5'd10};
		rom[ 602  ] = { 5'd0,	5'd6,	5'd6,	5'd7};
		rom[ 603  ] = { 5'd18,	5'd0,	5'd6,	5'd6};
		rom[ 604  ] = { 5'd3,	5'd1,	5'd18,	5'd3};
		rom[ 605  ] = { 5'd9,	5'd6,	5'd14,	5'd18};
		rom[ 606  ] = { 5'd0,	5'd0,	5'd6,	5'd6};
		rom[ 607  ] = { 5'd13,	5'd11,	5'd6,	5'd6};
		rom[ 608  ] = { 5'd0,	5'd20,	5'd24,	5'd3};
		rom[ 609  ] = { 5'd13,	5'd11,	5'd6,	5'd7};
		rom[ 610  ] = { 5'd4,	5'd12,	5'd10,	5'd6};
		rom[ 611  ] = { 5'd13,	5'd11,	5'd6,	5'd6};
		rom[ 612  ] = { 5'd5,	5'd11,	5'd6,	5'd7};
		rom[ 613  ] = { 5'd7,	5'd4,	5'd11,	5'd12};
		rom[ 614  ] = { 5'd6,	5'd15,	5'd10,	5'd4};
		rom[ 615  ] = { 5'd14,	5'd0,	5'd6,	5'd9};
		rom[ 616  ] = { 5'd4,	5'd0,	5'd6,	5'd9};
		rom[ 617  ] = { 5'd11,	5'd2,	5'd4,	5'd15};
		rom[ 618  ] = { 5'd0,	5'd0,	5'd20,	5'd3};
		rom[ 619  ] = { 5'd13,	5'd18,	5'd10,	5'd6};
		rom[ 620  ] = { 5'd2,	5'd7,	5'd6,	5'd11};
		rom[ 621  ] = { 5'd10,	5'd14,	5'd10,	5'd9};
		rom[ 622  ] = { 5'd8,	5'd2,	5'd4,	5'd9};
		rom[ 623  ] = { 5'd14,	5'd3,	5'd10,	5'd4};
		rom[ 624  ] = { 5'd6,	5'd6,	5'd12,	5'd6};
		rom[ 625  ] = { 5'd8,	5'd8,	5'd8,	5'd10};
		rom[ 626  ] = { 5'd7,	5'd4,	5'd4,	5'd16};
		rom[ 627  ] = { 5'd8,	5'd8,	5'd9,	5'd4};
		rom[ 628  ] = { 5'd5,	5'd2,	5'd14,	5'd9};
		rom[ 629  ] = { 5'd3,	5'd16,	5'd19,	5'd8};
		rom[ 630  ] = { 5'd0,	5'd0,	5'd10,	5'd8};
		rom[ 631  ] = { 5'd5,	5'd2,	5'd16,	5'd18};
		rom[ 632  ] = { 5'd0,	5'd11,	5'd24,	5'd11};
		rom[ 633  ] = { 5'd3,	5'd3,	5'd18,	5'd5};
		rom[ 634  ] = { 5'd1,	5'd16,	5'd18,	5'd3};
		rom[ 635  ] = { 5'd5,	5'd17,	5'd18,	5'd3};
		rom[ 636  ] = { 5'd1,	5'd13,	5'd9,	5'd6};
		rom[ 637  ] = { 5'd1,	5'd9,	5'd23,	5'd10};
		rom[ 638  ] = { 5'd3,	5'd7,	5'd18,	5'd3};
		rom[ 639  ] = { 5'd6,	5'd8,	5'd12,	5'd3};
		rom[ 640  ] = { 5'd6,	5'd2,	5'd3,	5'd22};
		rom[ 641  ] = { 5'd14,	5'd17,	5'd10,	5'd6};
		rom[ 642  ] = { 5'd1,	5'd18,	5'd10,	5'd6};
		rom[ 643  ] = { 5'd11,	5'd3,	5'd6,	5'd12};
		rom[ 644  ] = { 5'd10,	5'd6,	5'd4,	5'd9};
		rom[ 645  ] = { 5'd11,	5'd0,	5'd6,	5'd9};
		rom[ 646  ] = { 5'd7,	5'd0,	5'd6,	5'd9};
		rom[ 647  ] = { 5'd12,	5'd10,	5'd9,	5'd6};
		rom[ 648  ] = { 5'd2,	5'd11,	5'd6,	5'd9};
		rom[ 649  ] = { 5'd14,	5'd5,	5'd3,	5'd19};
		rom[ 650  ] = { 5'd6,	5'd6,	5'd9,	5'd6};
		rom[ 651  ] = { 5'd14,	5'd5,	5'd3,	5'd19};
		rom[ 652  ] = { 5'd0,	5'd3,	5'd6,	5'd9};
		rom[ 653  ] = { 5'd5,	5'd21,	5'd18,	5'd3};
		rom[ 654  ] = { 5'd1,	5'd10,	5'd18,	5'd4};
		rom[ 655  ] = { 5'd13,	5'd4,	5'd8,	5'd10};
		rom[ 656  ] = { 5'd7,	5'd8,	5'd9,	5'd6};
		rom[ 657  ] = { 5'd12,	5'd9,	5'd9,	5'd8};
		rom[ 658  ] = { 5'd0,	5'd6,	5'd5,	5'd12};
		rom[ 659  ] = { 5'd7,	5'd6,	5'd14,	5'd6};
		rom[ 660  ] = { 5'd7,	5'd5,	5'd3,	5'd19};
		rom[ 661  ] = { 5'd8,	5'd4,	5'd15,	5'd20};
		rom[ 662  ] = { 5'd1,	5'd4,	5'd15,	5'd20};
		rom[ 663  ] = { 5'd13,	5'd10,	5'd6,	5'd6};
		rom[ 664  ] = { 5'd5,	5'd10,	5'd6,	5'd6};
		rom[ 665  ] = { 5'd14,	5'd2,	5'd6,	5'd14};
		rom[ 666  ] = { 5'd4,	5'd2,	5'd6,	5'd14};
		rom[ 667  ] = { 5'd12,	5'd4,	5'd6,	5'd7};
		rom[ 668  ] = { 5'd9,	5'd4,	5'd6,	5'd9};
		rom[ 669  ] = { 5'd11,	5'd4,	5'd8,	5'd10};
		rom[ 670  ] = { 5'd5,	5'd4,	5'd8,	5'd10};
		rom[ 671  ] = { 5'd8,	5'd18,	5'd10,	5'd6};
		rom[ 672  ] = { 5'd1,	5'd18,	5'd21,	5'd6};
		rom[ 673  ] = { 5'd9,	5'd2,	5'd12,	5'd6};
		rom[ 674  ] = { 5'd3,	5'd2,	5'd12,	5'd6};
		rom[ 675  ] = { 5'd12,	5'd5,	5'd12,	5'd6};
		rom[ 676  ] = { 5'd8,	5'd8,	5'd6,	5'd9};
		rom[ 677  ] = { 5'd2,	5'd7,	5'd20,	5'd6};
		rom[ 678  ] = { 5'd0,	5'd5,	5'd12,	5'd6};
		rom[ 679  ] = { 5'd14,	5'd14,	5'd8,	5'd10};
		rom[ 680  ] = { 5'd2,	5'd14,	5'd8,	5'd10};
		rom[ 681  ] = { 5'd2,	5'd11,	5'd20,	5'd13};
		rom[ 682  ] = { 5'd6,	5'd9,	5'd12,	5'd5};
		rom[ 683  ] = { 5'd5,	5'd6,	5'd16,	5'd6};
		rom[ 684  ] = { 5'd1,	5'd19,	5'd9,	5'd4};
		rom[ 685  ] = { 5'd7,	5'd5,	5'd12,	5'd5};
		rom[ 686  ] = { 5'd3,	5'd5,	5'd14,	5'd12};
		rom[ 687  ] = { 5'd9,	5'd4,	5'd9,	5'd6};
		rom[ 688  ] = { 5'd2,	5'd6,	5'd19,	5'd3};
		rom[ 689  ] = { 5'd18,	5'd10,	5'd6,	5'd9};
		rom[ 690  ] = { 5'd3,	5'd7,	5'd18,	5'd2};
		rom[ 691  ] = { 5'd20,	5'd2,	5'd4,	5'd18};
		rom[ 692  ] = { 5'd2,	5'd18,	5'd20,	5'd3};
		rom[ 693  ] = { 5'd1,	5'd9,	5'd22,	5'd3};
		rom[ 694  ] = { 5'd0,	5'd2,	5'd4,	5'd18};
		rom[ 695  ] = { 5'd19,	5'd0,	5'd4,	5'd23};
		rom[ 696  ] = { 5'd0,	5'd3,	5'd6,	5'd19};
		rom[ 697  ] = { 5'd18,	5'd2,	5'd6,	5'd9};
		rom[ 698  ] = { 5'd0,	5'd5,	5'd10,	5'd6};
		rom[ 699  ] = { 5'd7,	5'd0,	5'd12,	5'd12};
		rom[ 700  ] = { 5'd0,	5'd3,	5'd24,	5'd6};
		rom[ 701  ] = { 5'd10,	5'd14,	5'd4,	5'd10};
		rom[ 702  ] = { 5'd8,	5'd9,	5'd4,	5'd15};
		rom[ 703  ] = { 5'd4,	5'd11,	5'd17,	5'd6};
		rom[ 704  ] = { 5'd2,	5'd5,	5'd18,	5'd8};
		rom[ 705  ] = { 5'd7,	5'd6,	5'd14,	5'd6};
		rom[ 706  ] = { 5'd3,	5'd6,	5'd14,	5'd6};
		rom[ 707  ] = { 5'd16,	5'd5,	5'd3,	5'd18};
		rom[ 708  ] = { 5'd5,	5'd5,	5'd3,	5'd18};
		rom[ 709  ] = { 5'd10,	5'd10,	5'd14,	5'd4};
		rom[ 710  ] = { 5'd4,	5'd10,	5'd9,	5'd4};
		rom[ 711  ] = { 5'd2,	5'd0,	5'd18,	5'd9};
		rom[ 712  ] = { 5'd6,	5'd3,	5'd12,	5'd8};
		rom[ 713  ] = { 5'd1,	5'd1,	5'd8,	5'd5};
		rom[ 714  ] = { 5'd12,	5'd7,	5'd7,	5'd8};
		rom[ 715  ] = { 5'd0,	5'd12,	5'd22,	5'd4};
		rom[ 716  ] = { 5'd15,	5'd6,	5'd4,	5'd15};
		rom[ 717  ] = { 5'd5,	5'd7,	5'd7,	5'd8};
		rom[ 718  ] = { 5'd8,	5'd18,	5'd9,	5'd4};
		rom[ 719  ] = { 5'd1,	5'd2,	5'd22,	5'd4};
		rom[ 720  ] = { 5'd17,	5'd3,	5'd6,	5'd17};
		rom[ 721  ] = { 5'd8,	5'd2,	5'd8,	5'd18};
		rom[ 722  ] = { 5'd17,	5'd0,	5'd6,	5'd12};
		rom[ 723  ] = { 5'd7,	5'd0,	5'd6,	5'd9};
		rom[ 724  ] = { 5'd15,	5'd5,	5'd9,	5'd12};
		rom[ 725  ] = { 5'd2,	5'd22,	5'd18,	5'd2};
		rom[ 726  ] = { 5'd10,	5'd10,	5'd12,	5'd6};
		rom[ 727  ] = { 5'd0,	5'd1,	5'd4,	5'd11};
		rom[ 728  ] = { 5'd20,	5'd0,	5'd4,	5'd10};
		rom[ 729  ] = { 5'd1,	5'd3,	5'd6,	5'd17};
		rom[ 730  ] = { 5'd15,	5'd15,	5'd9,	5'd6};
		rom[ 731  ] = { 5'd0,	5'd13,	5'd8,	5'd9};
		rom[ 732  ] = { 5'd16,	5'd8,	5'd6,	5'd12};
		rom[ 733  ] = { 5'd2,	5'd8,	5'd6,	5'd12};
		rom[ 734  ] = { 5'd10,	5'd2,	5'd4,	5'd15};
		rom[ 735  ] = { 5'd1,	5'd5,	5'd19,	5'd3};
		rom[ 736  ] = { 5'd11,	5'd8,	5'd9,	5'd7};
		rom[ 737  ] = { 5'd3,	5'd8,	5'd12,	5'd9};
		rom[ 738  ] = { 5'd3,	5'd6,	5'd18,	5'd3};
		rom[ 739  ] = { 5'd10,	5'd0,	5'd4,	5'd12};
		rom[ 740  ] = { 5'd3,	5'd9,	5'd18,	5'd14};
		rom[ 741  ] = { 5'd0,	5'd0,	5'd4,	5'd9};
		rom[ 742  ] = { 5'd12,	5'd5,	5'd4,	5'd18};
		rom[ 743  ] = { 5'd8,	5'd5,	5'd4,	5'd18};
		rom[ 744  ] = { 5'd10,	5'd5,	5'd6,	5'd10};
		rom[ 745  ] = { 5'd9,	5'd4,	5'd4,	5'd11};
		rom[ 746  ] = { 5'd4,	5'd16,	5'd18,	5'd3};
		rom[ 747  ] = { 5'd0,	5'd16,	5'd20,	5'd3};
		rom[ 748  ] = { 5'd9,	5'd9,	5'd6,	5'd12};
		rom[ 749  ] = { 5'd8,	5'd13,	5'd8,	5'd8};
		rom[ 750  ] = { 5'd13,	5'd10,	5'd3,	5'd12};
		rom[ 751  ] = { 5'd5,	5'd9,	5'd14,	5'd14};
		rom[ 752  ] = { 5'd0,	5'd0,	5'd24,	5'd10};
		rom[ 753  ] = { 5'd1,	5'd11,	5'd18,	5'd2};
		rom[ 754  ] = { 5'd19,	5'd5,	5'd5,	5'd12};
		rom[ 755  ] = { 5'd0,	5'd5,	5'd5,	5'd12};
		rom[ 756  ] = { 5'd16,	5'd6,	5'd8,	5'd18};
		rom[ 757  ] = { 5'd0,	5'd6,	5'd8,	5'd18};
		rom[ 758  ] = { 5'd12,	5'd5,	5'd12,	5'd12};
		rom[ 759  ] = { 5'd7,	5'd6,	5'd6,	5'd9};
		rom[ 760  ] = { 5'd9,	5'd13,	5'd6,	5'd11};
		rom[ 761  ] = { 5'd0,	5'd5,	5'd12,	5'd12};
		rom[ 762  ] = { 5'd1,	5'd2,	5'd23,	5'd3};
		rom[ 763  ] = { 5'd1,	5'd15,	5'd19,	5'd3};
		rom[ 764  ] = { 5'd13,	5'd17,	5'd11,	5'd4};
		rom[ 765  ] = { 5'd0,	5'd13,	5'd8,	5'd5};
		rom[ 766  ] = { 5'd12,	5'd10,	5'd10,	5'd4};
		rom[ 767  ] = { 5'd4,	5'd6,	5'd9,	5'd9};
		rom[ 768  ] = { 5'd15,	5'd14,	5'd9,	5'd6};
		rom[ 769  ] = { 5'd1,	5'd12,	5'd9,	5'd6};
		rom[ 770  ] = { 5'd3,	5'd10,	5'd20,	5'd8};
		rom[ 771  ] = { 5'd2,	5'd0,	5'd9,	5'd18};
		rom[ 772  ] = { 5'd13,	5'd11,	5'd9,	5'd10};
		rom[ 773  ] = { 5'd1,	5'd2,	5'd8,	5'd5};
		rom[ 774  ] = { 5'd3,	5'd4,	5'd21,	5'd6};
		rom[ 775  ] = { 5'd7,	5'd0,	5'd10,	5'd14};
		rom[ 776  ] = { 5'd12,	5'd17,	5'd12,	5'd4};
		rom[ 777  ] = { 5'd0,	5'd6,	5'd23,	5'd4};
		rom[ 778  ] = { 5'd13,	5'd10,	5'd8,	5'd10};
		rom[ 779  ] = { 5'd0,	5'd16,	5'd18,	5'd3};
		rom[ 780  ] = { 5'd15,	5'd16,	5'd9,	5'd4};
		rom[ 781  ] = { 5'd0,	5'd16,	5'd9,	5'd4};
		rom[ 782  ] = { 5'd13,	5'd11,	5'd6,	5'd6};
		rom[ 783  ] = { 5'd5,	5'd11,	5'd6,	5'd6};
		rom[ 784  ] = { 5'd0,	5'd3,	5'd24,	5'd6};
		rom[ 785  ] = { 5'd2,	5'd4,	5'd18,	5'd3};
		rom[ 786  ] = { 5'd0,	5'd0,	5'd24,	5'd4};
		rom[ 787  ] = { 5'd1,	5'd16,	5'd18,	5'd3};
		rom[ 788  ] = { 5'd15,	5'd15,	5'd9,	5'd6};
		rom[ 789  ] = { 5'd0,	5'd15,	5'd9,	5'd6};
		rom[ 790  ] = { 5'd6,	5'd17,	5'd18,	5'd3};
		rom[ 791  ] = { 5'd8,	5'd8,	5'd6,	5'd10};
		rom[ 792  ] = { 5'd10,	5'd6,	5'd6,	5'd9};
		rom[ 793  ] = { 5'd8,	5'd8,	5'd5,	5'd8};
		rom[ 794  ] = { 5'd12,	5'd8,	5'd6,	5'd8};
		rom[ 795  ] = { 5'd6,	5'd5,	5'd6,	5'd11};
		rom[ 796  ] = { 5'd13,	5'd6,	5'd8,	5'd9};
		rom[ 797  ] = { 5'd1,	5'd7,	5'd21,	5'd6};
		rom[ 798  ] = { 5'd15,	5'd5,	5'd3,	5'd12};
		rom[ 799  ] = { 5'd6,	5'd9,	5'd11,	5'd12};
		rom[ 800  ] = { 5'd13,	5'd8,	5'd10,	5'd8};
		rom[ 801  ] = { 5'd5,	5'd8,	5'd12,	5'd3};
		rom[ 802  ] = { 5'd6,	5'd11,	5'd18,	5'd4};
		rom[ 803  ] = { 5'd0,	5'd0,	5'd22,	5'd22};
		rom[ 804  ] = { 5'd11,	5'd2,	5'd6,	5'd8};
		rom[ 805  ] = { 5'd9,	5'd0,	5'd6,	5'd9};
		rom[ 806  ] = { 5'd10,	5'd0,	5'd6,	5'd9};
		rom[ 807  ] = { 5'd8,	5'd3,	5'd6,	5'd14};
		rom[ 808  ] = { 5'd3,	5'd10,	5'd18,	5'd8};
		rom[ 809  ] = { 5'd10,	5'd0,	5'd3,	5'd14};
		rom[ 810  ] = { 5'd4,	5'd3,	5'd16,	5'd20};
		rom[ 811  ] = { 5'd9,	5'd4,	5'd6,	5'd10};
		rom[ 812  ] = { 5'd5,	5'd0,	5'd16,	5'd4};
		rom[ 813  ] = { 5'd2,	5'd5,	5'd18,	5'd4};
		rom[ 814  ] = { 5'd13,	5'd0,	5'd6,	5'd9};
		rom[ 815  ] = { 5'd8,	5'd4,	5'd8,	5'd5};
		rom[ 816  ] = { 5'd12,	5'd10,	5'd10,	5'd4};
		rom[ 817  ] = { 5'd2,	5'd10,	5'd10,	5'd4};
		rom[ 818  ] = { 5'd7,	5'd11,	5'd12,	5'd5};
		rom[ 819  ] = { 5'd3,	5'd10,	5'd8,	5'd10};
		rom[ 820  ] = { 5'd11,	5'd12,	5'd9,	5'd8};
		rom[ 821  ] = { 5'd0,	5'd21,	5'd24,	5'd3};
		rom[ 822  ] = { 5'd3,	5'd20,	5'd18,	5'd4};
		rom[ 823  ] = { 5'd1,	5'd15,	5'd9,	5'd6};
		rom[ 824  ] = { 5'd11,	5'd17,	5'd10,	5'd4};
		rom[ 825  ] = { 5'd9,	5'd12,	5'd4,	5'd12};
		rom[ 826  ] = { 5'd9,	5'd6,	5'd9,	5'd6};
		rom[ 827  ] = { 5'd1,	5'd13,	5'd6,	5'd9};
		rom[ 828  ] = { 5'd6,	5'd16,	5'd12,	5'd4};
		rom[ 829  ] = { 5'd1,	5'd5,	5'd20,	5'd3};
		rom[ 830  ] = { 5'd8,	5'd1,	5'd9,	5'd9};
		rom[ 831  ] = { 5'd2,	5'd19,	5'd9,	5'd4};
		rom[ 832  ] = { 5'd11,	5'd1,	5'd4,	5'd18};
		rom[ 833  ] = { 5'd7,	5'd2,	5'd8,	5'd12};
		rom[ 834  ] = { 5'd11,	5'd10,	5'd9,	5'd8};
		rom[ 835  ] = { 5'd5,	5'd11,	5'd12,	5'd5};
		rom[ 836  ] = { 5'd11,	5'd9,	5'd9,	5'd6};
		rom[ 837  ] = { 5'd5,	5'd10,	5'd6,	5'd9};
		rom[ 838  ] = { 5'd4,	5'd7,	5'd5,	5'd12};
		rom[ 839  ] = { 5'd2,	5'd0,	5'd21,	5'd6};
		rom[ 840  ] = { 5'd7,	5'd6,	5'd10,	5'd6};
		rom[ 841  ] = { 5'd9,	5'd0,	5'd6,	5'd15};
		rom[ 842  ] = { 5'd2,	5'd2,	5'd18,	5'd2};
		rom[ 843  ] = { 5'd8,	5'd17,	5'd8,	5'd6};
		rom[ 844  ] = { 5'd3,	5'd0,	5'd18,	5'd2};
		rom[ 845  ] = { 5'd8,	5'd0,	5'd9,	5'd6};
		rom[ 846  ] = { 5'd0,	5'd17,	5'd18,	5'd3};
		rom[ 847  ] = { 5'd6,	5'd7,	5'd12,	5'd5};
		rom[ 848  ] = { 5'd0,	5'd3,	5'd6,	5'd9};
		rom[ 849  ] = { 5'd20,	5'd2,	5'd4,	5'd9};
		rom[ 850  ] = { 5'd0,	5'd2,	5'd4,	5'd9};
		rom[ 851  ] = { 5'd0,	5'd1,	5'd24,	5'd4};
		rom[ 852  ] = { 5'd0,	5'd16,	5'd9,	5'd6};
		rom[ 853  ] = { 5'd14,	5'd13,	5'd9,	5'd6};
		rom[ 854  ] = { 5'd0,	5'd15,	5'd19,	5'd3};
		rom[ 855  ] = { 5'd1,	5'd5,	5'd22,	5'd12};
		rom[ 856  ] = { 5'd5,	5'd13,	5'd6,	5'd6};
		rom[ 857  ] = { 5'd4,	5'd2,	5'd20,	5'd3};
		rom[ 858  ] = { 5'd8,	5'd14,	5'd6,	5'd10};
		rom[ 859  ] = { 5'd6,	5'd12,	5'd16,	5'd6};
		rom[ 860  ] = { 5'd2,	5'd13,	5'd8,	5'd9};
		rom[ 861  ] = { 5'd11,	5'd8,	5'd6,	5'd14};
		rom[ 862  ] = { 5'd2,	5'd12,	5'd16,	5'd6};
		rom[ 863  ] = { 5'd5,	5'd16,	5'd16,	5'd8};
		rom[ 864  ] = { 5'd9,	5'd1,	5'd4,	5'd12};
		rom[ 865  ] = { 5'd8,	5'd2,	5'd8,	5'd10};
		rom[ 866  ] = { 5'd6,	5'd6,	5'd12,	5'd6};
		rom[ 867  ] = { 5'd10,	5'd7,	5'd6,	5'd9};
		rom[ 868  ] = { 5'd0,	5'd0,	5'd8,	5'd12};
		rom[ 869  ] = { 5'd18,	5'd8,	5'd6,	5'd9};
		rom[ 870  ] = { 5'd2,	5'd12,	5'd6,	5'd6};
		rom[ 871  ] = { 5'd3,	5'd21,	5'd21,	5'd3};
		rom[ 872  ] = { 5'd2,	5'd0,	5'd16,	5'd6};
		rom[ 873  ] = { 5'd13,	5'd6,	5'd7,	5'd6};
		rom[ 874  ] = { 5'd6,	5'd4,	5'd4,	5'd14};
		rom[ 875  ] = { 5'd9,	5'd7,	5'd6,	5'd9};
		rom[ 876  ] = { 5'd7,	5'd8,	5'd6,	5'd14};
		rom[ 877  ] = { 5'd18,	5'd8,	5'd4,	5'd16};
		rom[ 878  ] = { 5'd9,	5'd14,	5'd6,	5'd10};
		rom[ 879  ] = { 5'd6,	5'd11,	5'd12,	5'd5};
		rom[ 880  ] = { 5'd0,	5'd12,	5'd23,	5'd3};
		rom[ 881  ] = { 5'd13,	5'd0,	5'd6,	5'd12};
		rom[ 882  ] = { 5'd0,	5'd10,	5'd12,	5'd5};
		rom[ 883  ] = { 5'd13,	5'd2,	5'd10,	5'd4};
		rom[ 884  ] = { 5'd5,	5'd0,	5'd6,	5'd12};
		rom[ 885  ] = { 5'd11,	5'd6,	5'd9,	5'd6};
		rom[ 886  ] = { 5'd4,	5'd6,	5'd9,	5'd6};
		rom[ 887  ] = { 5'd6,	5'd11,	5'd18,	5'd13};
		rom[ 888  ] = { 5'd0,	5'd11,	5'd18,	5'd13};
		rom[ 889  ] = { 5'd12,	5'd16,	5'd12,	5'd6};
		rom[ 890  ] = { 5'd0,	5'd6,	5'd21,	5'd3};
		rom[ 891  ] = { 5'd12,	5'd16,	5'd12,	5'd6};
		rom[ 892  ] = { 5'd5,	5'd7,	5'd6,	5'd14};
		rom[ 893  ] = { 5'd5,	5'd10,	5'd19,	5'd2};
		rom[ 894  ] = { 5'd5,	5'd4,	5'd14,	5'd4};
		rom[ 895  ] = { 5'd3,	5'd18,	5'd18,	5'd4};
		rom[ 896  ] = { 5'd7,	5'd0,	5'd4,	5'd9};
		rom[ 897  ] = { 5'd13,	5'd3,	5'd11,	5'd4};
		rom[ 898  ] = { 5'd2,	5'd0,	5'd9,	5'd6};
		rom[ 899  ] = { 5'd19,	5'd1,	5'd4,	5'd23};
		rom[ 900  ] = { 5'd1,	5'd1,	5'd4,	5'd23};
		rom[ 901  ] = { 5'd5,	5'd16,	5'd18,	5'd3};
		rom[ 902  ] = { 5'd0,	5'd3,	5'd11,	5'd4};
		rom[ 903  ] = { 5'd2,	5'd16,	5'd20,	5'd3};
		rom[ 904  ] = { 5'd5,	5'd3,	5'd13,	5'd4};
		rom[ 905  ] = { 5'd1,	5'd9,	5'd22,	5'd15};
		rom[ 906  ] = { 5'd3,	5'd4,	5'd14,	5'd3};
		rom[ 907  ] = { 5'd8,	5'd7,	5'd10,	5'd4};
		rom[ 908  ] = { 5'd6,	5'd7,	5'd10,	5'd4};
		rom[ 909  ] = { 5'd10,	5'd4,	5'd6,	5'd9};
		rom[ 910  ] = { 5'd1,	5'd12,	5'd9,	5'd6};
		rom[ 911  ] = { 5'd8,	5'd3,	5'd8,	5'd10};
		rom[ 912  ] = { 5'd3,	5'd6,	5'd16,	5'd6};
		rom[ 913  ] = { 5'd5,	5'd6,	5'd14,	5'd6};
		rom[ 914  ] = { 5'd4,	5'd3,	5'd9,	5'd6};
		rom[ 915  ] = { 5'd6,	5'd3,	5'd18,	5'd2};
		rom[ 916  ] = { 5'd7,	5'd6,	5'd9,	5'd6};
		rom[ 917  ] = { 5'd0,	5'd1,	5'd24,	5'd3};
		rom[ 918  ] = { 5'd0,	5'd17,	5'd10,	5'd6};
		rom[ 919  ] = { 5'd3,	5'd18,	5'd18,	5'd3};
		rom[ 920  ] = { 5'd2,	5'd5,	5'd6,	5'd16};
		rom[ 921  ] = { 5'd7,	5'd6,	5'd11,	5'd6};
		rom[ 922  ] = { 5'd5,	5'd2,	5'd12,	5'd22};
		rom[ 923  ] = { 5'd10,	5'd7,	5'd4,	5'd10};
		rom[ 924  ] = { 5'd9,	5'd0,	5'd4,	5'd18};
		rom[ 925  ] = { 5'd18,	5'd8,	5'd6,	5'd9};
		rom[ 926  ] = { 5'd4,	5'd7,	5'd15,	5'd10};
		rom[ 927  ] = { 5'd10,	5'd5,	5'd6,	5'd9};
		rom[ 928  ] = { 5'd9,	5'd9,	5'd6,	5'd10};
		rom[ 929  ] = { 5'd11,	5'd14,	5'd6,	5'd10};
		rom[ 930  ] = { 5'd7,	5'd14,	5'd6,	5'd10};
		rom[ 931  ] = { 5'd4,	5'd8,	5'd16,	5'd9};
		rom[ 932  ] = { 5'd2,	5'd11,	5'd20,	5'd3};
		rom[ 933  ] = { 5'd13,	5'd0,	5'd4,	5'd13};
		rom[ 934  ] = { 5'd7,	5'd0,	5'd4,	5'd13};
		rom[ 935  ] = { 5'd3,	5'd1,	5'd18,	5'd7};
		rom[ 936  ] = { 5'd1,	5'd11,	5'd6,	5'd9};
		rom[ 937  ] = { 5'd8,	5'd18,	5'd9,	5'd6};
		rom[ 938  ] = { 5'd3,	5'd9,	5'd15,	5'd6};
		rom[ 939  ] = { 5'd5,	5'd10,	5'd19,	5'd2};
		rom[ 940  ] = { 5'd8,	5'd6,	5'd7,	5'd16};
		rom[ 941  ] = { 5'd9,	5'd14,	5'd9,	5'd6};
		rom[ 942  ] = { 5'd0,	5'd7,	5'd8,	5'd12};
		rom[ 943  ] = { 5'd6,	5'd4,	5'd18,	5'd3};
		rom[ 944  ] = { 5'd0,	5'd16,	5'd12,	5'd6};
		rom[ 945  ] = { 5'd13,	5'd13,	5'd9,	5'd4};
		rom[ 946  ] = { 5'd5,	5'd8,	5'd14,	5'd14};
		rom[ 947  ] = { 5'd1,	5'd16,	5'd22,	5'd6};
		rom[ 948  ] = { 5'd9,	5'd0,	5'd6,	5'd9};
		rom[ 949  ] = { 5'd9,	5'd5,	5'd10,	5'd10};
		rom[ 950  ] = { 5'd5,	5'd5,	5'd10,	5'd10};
		rom[ 951  ] = { 5'd4,	5'd6,	5'd16,	5'd6};
		rom[ 952  ] = { 5'd0,	5'd7,	5'd6,	5'd9};
		rom[ 953  ] = { 5'd16,	5'd10,	5'd8,	5'd14};
		rom[ 954  ] = { 5'd9,	5'd12,	5'd6,	5'd12};
		rom[ 955  ] = { 5'd8,	5'd10,	5'd8,	5'd12};
		rom[ 956  ] = { 5'd8,	5'd0,	5'd4,	5'd9};
		rom[ 957  ] = { 5'd10,	5'd4,	5'd8,	5'd16};
		rom[ 958  ] = { 5'd7,	5'd10,	5'd10,	5'd6};
		rom[ 959  ] = { 5'd5,	5'd6,	5'd14,	5'd14};
		rom[ 960  ] = { 5'd2,	5'd11,	5'd20,	5'd2};
		rom[ 961  ] = { 5'd18,	5'd8,	5'd4,	5'd16};
		rom[ 962  ] = { 5'd1,	5'd11,	5'd12,	5'd10};
		rom[ 963  ] = { 5'd6,	5'd9,	5'd12,	5'd4};
		rom[ 964  ] = { 5'd9,	5'd12,	5'd6,	5'd7};
		rom[ 965  ] = { 5'd10,	5'd4,	5'd8,	5'd16};
		rom[ 966  ] = { 5'd6,	5'd4,	5'd8,	5'd16};
		rom[ 967  ] = { 5'd8,	5'd9,	5'd9,	5'd6};
		rom[ 968  ] = { 5'd1,	5'd5,	5'd16,	5'd12};
		rom[ 969  ] = { 5'd9,	5'd9,	5'd6,	5'd8};
		rom[ 970  ] = { 5'd6,	5'd0,	5'd3,	5'd18};
		rom[ 971  ] = { 5'd17,	5'd9,	5'd5,	5'd14};
		rom[ 972  ] = { 5'd2,	5'd9,	5'd5,	5'd14};
		rom[ 973  ] = { 5'd7,	5'd4,	5'd10,	5'd6};
		rom[ 974  ] = { 5'd1,	5'd3,	5'd23,	5'd18};
		rom[ 975  ] = { 5'd1,	5'd1,	5'd21,	5'd3};
		rom[ 976  ] = { 5'd9,	5'd6,	5'd6,	5'd9};
		rom[ 977  ] = { 5'd3,	5'd18,	5'd12,	5'd6};
		rom[ 978  ] = { 5'd16,	5'd8,	5'd8,	5'd16};
		rom[ 979  ] = { 5'd0,	5'd19,	5'd24,	5'd4};
		rom[ 980  ] = { 5'd16,	5'd8,	5'd8,	5'd16};
		rom[ 981  ] = { 5'd0,	5'd8,	5'd8,	5'd16};
		rom[ 982  ] = { 5'd8,	5'd12,	5'd8,	5'd10};
		rom[ 983  ] = { 5'd5,	5'd7,	5'd5,	5'd8};
		rom[ 984  ] = { 5'd4,	5'd1,	5'd19,	5'd2};
		rom[ 985  ] = { 5'd0,	5'd12,	5'd24,	5'd9};
		rom[ 986  ] = { 5'd6,	5'd0,	5'd13,	5'd8};
		rom[ 987  ] = { 5'd0,	5'd0,	5'd24,	5'd3};
		rom[ 988  ] = { 5'd20,	5'd3,	5'd4,	5'd11};
		rom[ 989  ] = { 5'd8,	5'd6,	5'd6,	5'd9};
		rom[ 990  ] = { 5'd6,	5'd11,	5'd12,	5'd8};
		rom[ 991  ] = { 5'd0,	5'd8,	5'd12,	5'd6};
		rom[ 992  ] = { 5'd6,	5'd17,	5'd18,	5'd3};
		rom[ 993  ] = { 5'd0,	5'd14,	5'd9,	5'd6};
		rom[ 994  ] = { 5'd20,	5'd3,	5'd4,	5'd9};
		rom[ 995  ] = { 5'd0,	5'd3,	5'd4,	5'd9};
		rom[ 996  ] = { 5'd15,	5'd0,	5'd9,	5'd19};
		rom[ 997  ] = { 5'd0,	5'd0,	5'd9,	5'd19};
		rom[ 998  ] = { 5'd13,	5'd11,	5'd6,	5'd8};
		rom[ 999  ] = { 5'd5,	5'd11,	5'd6,	5'd8};
		rom[ 1000 ] = { 5'd5,	5'd11,	5'd19,	5'd3};
		rom[ 1001 ] = { 5'd3,	5'd20,	5'd18,	5'd4};
		rom[ 1002 ] = { 5'd6,	5'd6,	5'd16,	5'd6};
		rom[ 1003 ] = { 5'd6,	5'd0,	5'd9,	5'd6};
		rom[ 1004 ] = { 5'd10,	5'd3,	5'd4,	5'd14};
		rom[ 1005 ] = { 5'd1,	5'd5,	5'd15,	5'd12};
		rom[ 1006 ] = { 5'd11,	5'd12,	5'd8,	5'd5};
		rom[ 1007 ] = { 5'd5,	5'd0,	5'd6,	5'd9};
		rom[ 1008 ] = { 5'd12,	5'd0,	5'd6,	5'd9};
		rom[ 1009 ] = { 5'd5,	5'd5,	5'd12,	5'd8};
		rom[ 1010 ] = { 5'd13,	5'd12,	5'd11,	5'd6};
		rom[ 1011 ] = { 5'd0,	5'd13,	5'd21,	5'd3};
		rom[ 1012 ] = { 5'd8,	5'd1,	5'd8,	5'd12};
		rom[ 1013 ] = { 5'd1,	5'd0,	5'd6,	5'd12};
		rom[ 1014 ] = { 5'd2,	5'd2,	5'd21,	5'd2};
		rom[ 1015 ] = { 5'd2,	5'd2,	5'd19,	5'd3};
		rom[ 1016 ] = { 5'd17,	5'd10,	5'd6,	5'd14};
		rom[ 1017 ] = { 5'd1,	5'd10,	5'd6,	5'd14};
		rom[ 1018 ] = { 5'd7,	5'd6,	5'd14,	5'd14};
		rom[ 1019 ] = { 5'd0,	5'd12,	5'd9,	5'd6};
		rom[ 1020 ] = { 5'd15,	5'd14,	5'd8,	5'd9};
		rom[ 1021 ] = { 5'd1,	5'd1,	5'd22,	5'd4};
		rom[ 1022 ] = { 5'd9,	5'd11,	5'd9,	5'd6};
		rom[ 1023 ] = { 5'd0,	5'd15,	5'd18,	5'd3};
		rom[ 1024 ] = { 5'd16,	5'd14,	5'd7,	5'd9};
		rom[ 1025 ] = { 5'd4,	5'd3,	5'd16,	5'd4};
		rom[ 1026 ] = { 5'd7,	5'd6,	5'd12,	5'd5};
		rom[ 1027 ] = { 5'd9,	5'd6,	5'd4,	5'd9};
		rom[ 1028 ] = { 5'd12,	5'd1,	5'd4,	5'd10};
		rom[ 1029 ] = { 5'd8,	5'd1,	5'd4,	5'd10};
		rom[ 1030 ] = { 5'd15,	5'd15,	5'd6,	5'd9};
		rom[ 1031 ] = { 5'd3,	5'd15,	5'd6,	5'd9};
		rom[ 1032 ] = { 5'd15,	5'd1,	5'd3,	5'd19};
		rom[ 1033 ] = { 5'd1,	5'd3,	5'd6,	5'd9};
		rom[ 1034 ] = { 5'd15,	5'd0,	5'd3,	5'd19};
		rom[ 1035 ] = { 5'd6,	5'd3,	5'd12,	5'd4};
		rom[ 1036 ] = { 5'd10,	5'd5,	5'd4,	5'd9};
		rom[ 1037 ] = { 5'd6,	5'd0,	5'd3,	5'd19};
		rom[ 1038 ] = { 5'd11,	5'd1,	5'd3,	5'd12};
		rom[ 1039 ] = { 5'd6,	5'd7,	5'd10,	5'd5};
		rom[ 1040 ] = { 5'd11,	5'd3,	5'd3,	5'd18};
		rom[ 1041 ] = { 5'd9,	5'd3,	5'd6,	5'd12};
		rom[ 1042 ] = { 5'd3,	5'd7,	5'd19,	5'd3};
		rom[ 1043 ] = { 5'd2,	5'd7,	5'd18,	5'd3};
		rom[ 1044 ] = { 5'd3,	5'd13,	5'd18,	5'd4};
		rom[ 1045 ] = { 5'd3,	5'd5,	5'd6,	5'd9};
		rom[ 1046 ] = { 5'd4,	5'd1,	5'd20,	5'd4};
		rom[ 1047 ] = { 5'd0,	5'd1,	5'd20,	5'd4};
		rom[ 1048 ] = { 5'd10,	5'd15,	5'd6,	5'd6};
		rom[ 1049 ] = { 5'd0,	5'd2,	5'd24,	5'd8};
		rom[ 1050 ] = { 5'd5,	5'd5,	5'd18,	5'd3};
		rom[ 1051 ] = { 5'd8,	5'd15,	5'd6,	5'd6};
		rom[ 1052 ] = { 5'd11,	5'd12,	5'd8,	5'd5};
		rom[ 1053 ] = { 5'd5,	5'd12,	5'd8,	5'd5};
		rom[ 1054 ] = { 5'd5,	5'd0,	5'd14,	5'd6};
		rom[ 1055 ] = { 5'd10,	5'd2,	5'd4,	5'd15};
		rom[ 1056 ] = { 5'd10,	5'd7,	5'd5,	5'd12};
		rom[ 1057 ] = { 5'd7,	5'd9,	5'd8,	5'd14};
		rom[ 1058 ] = { 5'd1,	5'd5,	5'd22,	5'd6};
		rom[ 1059 ] = { 5'd0,	5'd5,	5'd6,	5'd6};
		rom[ 1060 ] = { 5'd12,	5'd17,	5'd9,	5'd4};
		rom[ 1061 ] = { 5'd2,	5'd18,	5'd19,	5'd3};
		rom[ 1062 ] = { 5'd12,	5'd17,	5'd9,	5'd4};
		rom[ 1063 ] = { 5'd1,	5'd17,	5'd18,	5'd3};
		rom[ 1064 ] = { 5'd12,	5'd17,	5'd9,	5'd4};
		rom[ 1065 ] = { 5'd0,	5'd0,	5'd24,	5'd3};
		rom[ 1066 ] = { 5'd5,	5'd0,	5'd14,	5'd4};
		rom[ 1067 ] = { 5'd6,	5'd14,	5'd9,	5'd6};
		rom[ 1068 ] = { 5'd14,	5'd13,	5'd6,	5'd9};
		rom[ 1069 ] = { 5'd5,	5'd20,	5'd13,	5'd4};
		rom[ 1070 ] = { 5'd9,	5'd9,	5'd6,	5'd12};
		rom[ 1071 ] = { 5'd1,	5'd10,	5'd21,	5'd3};
		rom[ 1072 ] = { 5'd8,	5'd8,	5'd9,	5'd6};
		rom[ 1073 ] = { 5'd3,	5'd10,	5'd9,	5'd7};
		rom[ 1074 ] = { 5'd12,	5'd10,	5'd10,	5'd8};
		rom[ 1075 ] = { 5'd0,	5'd15,	5'd24,	5'd3};
		rom[ 1076 ] = { 5'd8,	5'd5,	5'd9,	5'd6};
		rom[ 1077 ] = { 5'd4,	5'd13,	5'd6,	5'd9};
		rom[ 1078 ] = { 5'd12,	5'd17,	5'd9,	5'd4};
		rom[ 1079 ] = { 5'd9,	5'd12,	5'd6,	5'd6};
		rom[ 1080 ] = { 5'd9,	5'd9,	5'd14,	5'd10};
		rom[ 1081 ] = { 5'd1,	5'd9,	5'd14,	5'd10};
		rom[ 1082 ] = { 5'd8,	5'd7,	5'd9,	5'd17};
		rom[ 1083 ] = { 5'd3,	5'd4,	5'd6,	5'd20};
		rom[ 1084 ] = { 5'd7,	5'd8,	5'd10,	5'd4};
		rom[ 1085 ] = { 5'd10,	5'd7,	5'd4,	5'd9};
		rom[ 1086 ] = { 5'd10,	5'd15,	5'd6,	5'd9};
		rom[ 1087 ] = { 5'd3,	5'd8,	5'd6,	5'd16};
		rom[ 1088 ] = { 5'd12,	5'd17,	5'd9,	5'd4};
		rom[ 1089 ] = { 5'd3,	5'd17,	5'd9,	5'd4};
		rom[ 1090 ] = { 5'd10,	5'd1,	5'd9,	5'd6};
		rom[ 1091 ] = { 5'd5,	5'd7,	5'd4,	5'd10};
		rom[ 1092 ] = { 5'd7,	5'd5,	5'd12,	5'd6};
		rom[ 1093 ] = { 5'd6,	5'd4,	5'd9,	5'd8};
		rom[ 1094 ] = { 5'd12,	5'd16,	5'd10,	5'd8};
		rom[ 1095 ] = { 5'd2,	5'd16,	5'd10,	5'd8};
		rom[ 1096 ] = { 5'd0,	5'd0,	5'd24,	5'd4};
		rom[ 1097 ] = { 5'd0,	5'd6,	5'd9,	5'd6};
		rom[ 1098 ] = { 5'd0,	5'd4,	5'd24,	5'd6};
		rom[ 1099 ] = { 5'd5,	5'd0,	5'd11,	5'd4};
		rom[ 1100 ] = { 5'd1,	5'd1,	5'd22,	5'd4};
		rom[ 1101 ] = { 5'd9,	5'd6,	5'd6,	5'd18};
		rom[ 1102 ] = { 5'd2,	5'd9,	5'd20,	5'd4};
		rom[ 1103 ] = { 5'd5,	5'd2,	5'd14,	5'd14};
		rom[ 1104 ] = { 5'd4,	5'd2,	5'd16,	5'd6};
		rom[ 1105 ] = { 5'd2,	5'd3,	5'd19,	5'd3};
		rom[ 1106 ] = { 5'd7,	5'd1,	5'd10,	5'd4};
		rom[ 1107 ] = { 5'd0,	5'd9,	5'd4,	5'd15};
		rom[ 1108 ] = { 5'd2,	5'd10,	5'd21,	5'd3};
		rom[ 1109 ] = { 5'd3,	5'd0,	5'd6,	5'd6};
		rom[ 1110 ] = { 5'd6,	5'd4,	5'd14,	5'd9};
		rom[ 1111 ] = { 5'd9,	5'd1,	5'd6,	5'd9};
		rom[ 1112 ] = { 5'd15,	5'd8,	5'd9,	5'd9};
		rom[ 1113 ] = { 5'd8,	5'd0,	5'd4,	5'd21};
		rom[ 1114 ] = { 5'd3,	5'd22,	5'd19,	5'd2};
		rom[ 1115 ] = { 5'd2,	5'd15,	5'd20,	5'd3};
		rom[ 1116 ] = { 5'd19,	5'd0,	5'd4,	5'd13};
		rom[ 1117 ] = { 5'd1,	5'd7,	5'd8,	5'd8};
		rom[ 1118 ] = { 5'd14,	5'd14,	5'd6,	5'd9};
		rom[ 1119 ] = { 5'd4,	5'd14,	5'd6,	5'd9};
		rom[ 1120 ] = { 5'd14,	5'd5,	5'd4,	5'd10};
		rom[ 1121 ] = { 5'd6,	5'd5,	5'd4,	5'd10};
		rom[ 1122 ] = { 5'd14,	5'd5,	5'd6,	5'd6};
		rom[ 1123 ] = { 5'd4,	5'd5,	5'd6,	5'd6};
		rom[ 1124 ] = { 5'd0,	5'd2,	5'd24,	5'd21};
		rom[ 1125 ] = { 5'd1,	5'd2,	5'd6,	5'd13};
		rom[ 1126 ] = { 5'd20,	5'd0,	5'd4,	5'd21};
		rom[ 1127 ] = { 5'd0,	5'd4,	5'd4,	5'd20};
		rom[ 1128 ] = { 5'd8,	5'd16,	5'd9,	5'd6};
		rom[ 1129 ] = { 5'd7,	5'd0,	5'd6,	5'd9};
		rom[ 1130 ] = { 5'd16,	5'd12,	5'd7,	5'd9};
		rom[ 1131 ] = { 5'd5,	5'd21,	5'd14,	5'd3};
		rom[ 1132 ] = { 5'd11,	5'd5,	5'd6,	5'd9};
		rom[ 1133 ] = { 5'd10,	5'd5,	5'd4,	5'd10};
		rom[ 1134 ] = { 5'd10,	5'd6,	5'd6,	5'd9};
		rom[ 1135 ] = { 5'd7,	5'd5,	5'd6,	5'd9};
		rom[ 1136 ] = { 5'd14,	5'd14,	5'd10,	5'd4};
		rom[ 1137 ] = { 5'd5,	5'd5,	5'd14,	5'd14};
		rom[ 1138 ] = { 5'd12,	5'd8,	5'd12,	5'd6};
		rom[ 1139 ] = { 5'd6,	5'd6,	5'd12,	5'd12};
		rom[ 1140 ] = { 5'd11,	5'd13,	5'd6,	5'd10};
		rom[ 1141 ] = { 5'd1,	5'd10,	5'd20,	5'd8};
		rom[ 1142 ] = { 5'd15,	5'd13,	5'd9,	5'd6};
		rom[ 1143 ] = { 5'd9,	5'd0,	5'd6,	5'd9};
		rom[ 1144 ] = { 5'd10,	5'd1,	5'd5,	5'd14};
		rom[ 1145 ] = { 5'd3,	5'd4,	5'd16,	5'd6};
		rom[ 1146 ] = { 5'd16,	5'd3,	5'd8,	5'd9};
		rom[ 1147 ] = { 5'd7,	5'd13,	5'd6,	5'd10};
		rom[ 1148 ] = { 5'd15,	5'd13,	5'd9,	5'd6};
		rom[ 1149 ] = { 5'd0,	5'd13,	5'd9,	5'd6};
		rom[ 1150 ] = { 5'd13,	5'd16,	5'd9,	5'd6};
		rom[ 1151 ] = { 5'd2,	5'd16,	5'd9,	5'd6};
		rom[ 1152 ] = { 5'd5,	5'd16,	5'd18,	5'd3};
		rom[ 1153 ] = { 5'd1,	5'd16,	5'd18,	5'd3};
		rom[ 1154 ] = { 5'd5,	5'd0,	5'd18,	5'd3};
		rom[ 1155 ] = { 5'd1,	5'd1,	5'd19,	5'd2};
		rom[ 1156 ] = { 5'd14,	5'd2,	5'd6,	5'd11};
		rom[ 1157 ] = { 5'd4,	5'd15,	5'd15,	5'd6};
		rom[ 1158 ] = { 5'd14,	5'd2,	5'd6,	5'd11};
		rom[ 1159 ] = { 5'd4,	5'd2,	5'd6,	5'd11};
		rom[ 1160 ] = { 5'd18,	5'd2,	5'd6,	5'd9};
		rom[ 1161 ] = { 5'd1,	5'd2,	5'd22,	5'd4};
		rom[ 1162 ] = { 5'd2,	5'd0,	5'd21,	5'd12};
		rom[ 1163 ] = { 5'd0,	5'd12,	5'd18,	5'd3};
		rom[ 1164 ] = { 5'd12,	5'd2,	5'd6,	5'd9};
		rom[ 1165 ] = { 5'd3,	5'd10,	5'd18,	5'd3};
		rom[ 1166 ] = { 5'd16,	5'd3,	5'd8,	5'd9};
		rom[ 1167 ] = { 5'd3,	5'd7,	5'd18,	5'd3};
		rom[ 1168 ] = { 5'd9,	5'd11,	5'd6,	5'd9};
		rom[ 1169 ] = { 5'd9,	5'd8,	5'd6,	5'd9};
		rom[ 1170 ] = { 5'd15,	5'd0,	5'd2,	5'd18};
		rom[ 1171 ] = { 5'd7,	5'd0,	5'd2,	5'd18};
		rom[ 1172 ] = { 5'd17,	5'd3,	5'd7,	5'd9};
		rom[ 1173 ] = { 5'd3,	5'd18,	5'd9,	5'd6};
		rom[ 1174 ] = { 5'd3,	5'd18,	5'd21,	5'd3};
		rom[ 1175 ] = { 5'd0,	5'd3,	5'd7,	5'd9};
		rom[ 1176 ] = { 5'd2,	5'd7,	5'd22,	5'd3};
		rom[ 1177 ] = { 5'd0,	5'd3,	5'd24,	5'd16};
		rom[ 1178 ] = { 5'd13,	5'd17,	5'd9,	5'd4};
		rom[ 1179 ] = { 5'd5,	5'd5,	5'd12,	5'd8};
		rom[ 1180 ] = { 5'd5,	5'd6,	5'd14,	5'd6};
		rom[ 1181 ] = { 5'd5,	5'd16,	5'd14,	5'd6};
		rom[ 1182 ] = { 5'd18,	5'd2,	5'd6,	5'd9};
		rom[ 1183 ] = { 5'd0,	5'd2,	5'd6,	5'd9};
		rom[ 1184 ] = { 5'd3,	5'd4,	5'd20,	5'd10};
		rom[ 1185 ] = { 5'd2,	5'd13,	5'd9,	5'd8};
		rom[ 1186 ] = { 5'd2,	5'd1,	5'd21,	5'd15};
		rom[ 1187 ] = { 5'd5,	5'd12,	5'd14,	5'd8};
		rom[ 1188 ] = { 5'd6,	5'd7,	5'd12,	5'd4};
		rom[ 1189 ] = { 5'd6,	5'd5,	5'd9,	5'd6};
		rom[ 1190 ] = { 5'd13,	5'd11,	5'd6,	5'd6};
		rom[ 1191 ] = { 5'd5,	5'd11,	5'd6,	5'd6};
		rom[ 1192 ] = { 5'd6,	5'd4,	5'd18,	5'd2};
		rom[ 1193 ] = { 5'd0,	5'd2,	5'd6,	5'd11};
		rom[ 1194 ] = { 5'd18,	5'd0,	5'd6,	5'd15};
		rom[ 1195 ] = { 5'd0,	5'd0,	5'd6,	5'd13};
		rom[ 1196 ] = { 5'd12,	5'd0,	5'd6,	5'd9};
		rom[ 1197 ] = { 5'd6,	5'd0,	5'd6,	5'd9};
		rom[ 1198 ] = { 5'd0,	5'd2,	5'd24,	5'd4};
		rom[ 1199 ] = { 5'd3,	5'd13,	5'd18,	5'd4};
		rom[ 1200 ] = { 5'd9,	5'd7,	5'd10,	5'd4};
		rom[ 1201 ] = { 5'd5,	5'd8,	5'd12,	5'd3};
		rom[ 1202 ] = { 5'd4,	5'd14,	5'd19,	5'd3};
		rom[ 1203 ] = { 5'd10,	5'd0,	5'd4,	5'd20};
		rom[ 1204 ] = { 5'd8,	5'd15,	5'd9,	5'd6};
		rom[ 1205 ] = { 5'd2,	5'd9,	5'd15,	5'd4};
		rom[ 1206 ] = { 5'd8,	5'd4,	5'd12,	5'd7};
		rom[ 1207 ] = { 5'd0,	5'd10,	5'd6,	5'd9};
		rom[ 1208 ] = { 5'd18,	5'd5,	5'd6,	5'd9};
		rom[ 1209 ] = { 5'd0,	5'd18,	5'd16,	5'd6};
		rom[ 1210 ] = { 5'd9,	5'd18,	5'd14,	5'd6};
		rom[ 1211 ] = { 5'd1,	5'd20,	5'd20,	5'd4};
		rom[ 1212 ] = { 5'd2,	5'd8,	5'd20,	5'd6};
		rom[ 1213 ] = { 5'd7,	5'd8,	5'd6,	5'd9};
		rom[ 1214 ] = { 5'd8,	5'd5,	5'd12,	5'd8};
		rom[ 1215 ] = { 5'd4,	5'd5,	5'd12,	5'd8};
		rom[ 1216 ] = { 5'd10,	5'd6,	5'd6,	5'd9};
		rom[ 1217 ] = { 5'd2,	5'd0,	5'd6,	5'd16};
		rom[ 1218 ] = { 5'd15,	5'd4,	5'd6,	5'd12};
		rom[ 1219 ] = { 5'd3,	5'd4,	5'd6,	5'd12};
		rom[ 1220 ] = { 5'd15,	5'd12,	5'd9,	5'd6};
		rom[ 1221 ] = { 5'd4,	5'd0,	5'd15,	5'd22};
		rom[ 1222 ] = { 5'd15,	5'd12,	5'd9,	5'd6};
		rom[ 1223 ] = { 5'd0,	5'd12,	5'd9,	5'd6};
		rom[ 1224 ] = { 5'd15,	5'd15,	5'd9,	5'd6};
		rom[ 1225 ] = { 5'd0,	5'd15,	5'd9,	5'd6};
		rom[ 1226 ] = { 5'd10,	5'd0,	5'd8,	5'd10};
		rom[ 1227 ] = { 5'd1,	5'd0,	5'd4,	5'd16};
		rom[ 1228 ] = { 5'd7,	5'd6,	5'd10,	5'd6};
		rom[ 1229 ] = { 5'd10,	5'd12,	5'd4,	5'd10};
		rom[ 1230 ] = { 5'd8,	5'd4,	5'd10,	5'd6};
		rom[ 1231 ] = { 5'd3,	5'd22,	5'd18,	5'd2};
		rom[ 1232 ] = { 5'd7,	5'd7,	5'd11,	5'd6};
		rom[ 1233 ] = { 5'd0,	5'd0,	5'd12,	5'd10};
		rom[ 1234 ] = { 5'd10,	5'd1,	5'd12,	5'd6};
		rom[ 1235 ] = { 5'd7,	5'd16,	5'd9,	5'd4};
		rom[ 1236 ] = { 5'd5,	5'd7,	5'd15,	5'd16};
		rom[ 1237 ] = { 5'd5,	5'd10,	5'd12,	5'd13};
		rom[ 1238 ] = { 5'd6,	5'd2,	5'd12,	5'd6};
		rom[ 1239 ] = { 5'd3,	5'd9,	5'd12,	5'd9};
		rom[ 1240 ] = { 5'd16,	5'd2,	5'd8,	5'd6};
		rom[ 1241 ] = { 5'd0,	5'd2,	5'd8,	5'd6};
		rom[ 1242 ] = { 5'd0,	5'd3,	5'd24,	5'd11};
		rom[ 1243 ] = { 5'd0,	5'd13,	5'd8,	5'd10};
		rom[ 1244 ] = { 5'd10,	5'd14,	5'd4,	5'd10};
		rom[ 1245 ] = { 5'd10,	5'd2,	5'd4,	5'd21};
		rom[ 1246 ] = { 5'd4,	5'd4,	5'd15,	5'd9};
		rom[ 1247 ] = { 5'd0,	5'd1,	5'd24,	5'd6};
		rom[ 1248 ] = { 5'd9,	5'd6,	5'd5,	5'd16};
		rom[ 1249 ] = { 5'd3,	5'd21,	5'd18,	5'd3};
		rom[ 1250 ] = { 5'd6,	5'd5,	5'd3,	5'd12};
		rom[ 1251 ] = { 5'd11,	5'd6,	5'd4,	5'd9};
		rom[ 1252 ] = { 5'd5,	5'd6,	5'd9,	5'd8};
		rom[ 1253 ] = { 5'd4,	5'd3,	5'd20,	5'd2};
		rom[ 1254 ] = { 5'd2,	5'd10,	5'd18,	5'd3};
		rom[ 1255 ] = { 5'd7,	5'd15,	5'd10,	5'd6};
		rom[ 1256 ] = { 5'd1,	5'd4,	5'd4,	5'd18};
		rom[ 1257 ] = { 5'd13,	5'd0,	5'd6,	5'd9};
		rom[ 1258 ] = { 5'd5,	5'd0,	5'd6,	5'd9};
		rom[ 1259 ] = { 5'd11,	5'd0,	5'd6,	5'd9};
		rom[ 1260 ] = { 5'd6,	5'd7,	5'd9,	5'd6};
		rom[ 1261 ] = { 5'd3,	5'd0,	5'd18,	5'd2};
		rom[ 1262 ] = { 5'd0,	5'd10,	5'd20,	5'd4};
		rom[ 1263 ] = { 5'd10,	5'd2,	5'd4,	5'd12};
		rom[ 1264 ] = { 5'd6,	5'd5,	5'd6,	5'd12};
		rom[ 1265 ] = { 5'd6,	5'd0,	5'd18,	5'd22};
		rom[ 1266 ] = { 5'd0,	5'd0,	5'd18,	5'd22};
		rom[ 1267 ] = { 5'd18,	5'd2,	5'd6,	5'd11};
		rom[ 1268 ] = { 5'd0,	5'd2,	5'd6,	5'd11};
		rom[ 1269 ] = { 5'd11,	5'd0,	5'd6,	5'd9};
		rom[ 1270 ] = { 5'd0,	5'd0,	5'd20,	5'd3};
		rom[ 1271 ] = { 5'd2,	5'd2,	5'd20,	5'd2};
		rom[ 1272 ] = { 5'd1,	5'd10,	5'd18,	5'd2};
		rom[ 1273 ] = { 5'd18,	5'd7,	5'd6,	5'd9};
		rom[ 1274 ] = { 5'd0,	5'd0,	5'd22,	5'd9};
		rom[ 1275 ] = { 5'd17,	5'd3,	5'd6,	5'd9};
		rom[ 1276 ] = { 5'd0,	5'd7,	5'd6,	5'd9};
		rom[ 1277 ] = { 5'd0,	5'd6,	5'd24,	5'd6};
		rom[ 1278 ] = { 5'd0,	5'd2,	5'd6,	5'd10};
		rom[ 1279 ] = { 5'd10,	5'd6,	5'd6,	5'd9};
		rom[ 1280 ] = { 5'd7,	5'd0,	5'd6,	5'd9};
		rom[ 1281 ] = { 5'd15,	5'd0,	5'd6,	5'd9};
		rom[ 1282 ] = { 5'd3,	5'd0,	5'd6,	5'd9};
		rom[ 1283 ] = { 5'd15,	5'd17,	5'd9,	5'd6};
		rom[ 1284 ] = { 5'd0,	5'd17,	5'd18,	5'd3};
		rom[ 1285 ] = { 5'd15,	5'd14,	5'd9,	5'd6};
		rom[ 1286 ] = { 5'd0,	5'd15,	5'd23,	5'd6};
		rom[ 1287 ] = { 5'd5,	5'd15,	5'd18,	5'd3};
		rom[ 1288 ] = { 5'd0,	5'd14,	5'd9,	5'd6};
		rom[ 1289 ] = { 5'd9,	5'd8,	5'd8,	5'd10};
		rom[ 1290 ] = { 5'd3,	5'd7,	5'd15,	5'd6};
		rom[ 1291 ] = { 5'd9,	5'd8,	5'd8,	5'd10};
		rom[ 1292 ] = { 5'd5,	5'd0,	5'd6,	5'd12};
		rom[ 1293 ] = { 5'd9,	5'd8,	5'd8,	5'd10};
		rom[ 1294 ] = { 5'd8,	5'd5,	5'd6,	5'd9};
		rom[ 1295 ] = { 5'd10,	5'd6,	5'd4,	5'd18};
		rom[ 1296 ] = { 5'd5,	5'd7,	5'd12,	5'd4};
		rom[ 1297 ] = { 5'd9,	5'd8,	5'd8,	5'd10};
		rom[ 1298 ] = { 5'd7,	5'd8,	5'd8,	5'd10};
		rom[ 1299 ] = { 5'd11,	5'd10,	5'd6,	5'd14};
		rom[ 1300 ] = { 5'd9,	5'd5,	5'd6,	5'd19};
		rom[ 1301 ] = { 5'd6,	5'd12,	5'd12,	5'd6};
		rom[ 1302 ] = { 5'd1,	5'd9,	5'd18,	5'd6};
		rom[ 1303 ] = { 5'd16,	5'd14,	5'd8,	5'd10};
		rom[ 1304 ] = { 5'd0,	5'd9,	5'd22,	5'd8};
		rom[ 1305 ] = { 5'd8,	5'd18,	5'd12,	5'd6};
		rom[ 1306 ] = { 5'd0,	5'd6,	5'd20,	5'd18};
		rom[ 1307 ] = { 5'd3,	5'd6,	5'd20,	5'd12};
		rom[ 1308 ] = { 5'd0,	5'd16,	5'd10,	5'd8};
		rom[ 1309 ] = { 5'd6,	5'd16,	5'd18,	5'd3};
		rom[ 1310 ] = { 5'd0,	5'd11,	5'd19,	5'd3};
		rom[ 1311 ] = { 5'd14,	5'd6,	5'd6,	5'd9};
		rom[ 1312 ] = { 5'd1,	5'd7,	5'd22,	5'd4};
		rom[ 1313 ] = { 5'd13,	5'd6,	5'd7,	5'd12};
		rom[ 1314 ] = { 5'd4,	5'd7,	5'd11,	5'd9};
		rom[ 1315 ] = { 5'd12,	5'd10,	5'd10,	5'd8};
		rom[ 1316 ] = { 5'd2,	5'd12,	5'd9,	5'd7};
		rom[ 1317 ] = { 5'd16,	5'd14,	5'd6,	5'd9};
		rom[ 1318 ] = { 5'd3,	5'd12,	5'd6,	5'd12};
		rom[ 1319 ] = { 5'd14,	5'd13,	5'd6,	5'd6};
		rom[ 1320 ] = { 5'd8,	5'd0,	5'd6,	5'd9};
		rom[ 1321 ] = { 5'd9,	5'd1,	5'd6,	5'd23};
		rom[ 1322 ] = { 5'd0,	5'd16,	5'd9,	5'd6};
		rom[ 1323 ] = { 5'd4,	5'd17,	5'd18,	5'd3};
		rom[ 1324 ] = { 5'd5,	5'd2,	5'd13,	5'd14};
		rom[ 1325 ] = { 5'd15,	5'd0,	5'd8,	5'd12};
		rom[ 1326 ] = { 5'd0,	5'd0,	5'd8,	5'd12};
		rom[ 1327 ] = { 5'd8,	5'd2,	5'd8,	5'd7};
		rom[ 1328 ] = { 5'd1,	5'd1,	5'd6,	5'd9};
		rom[ 1329 ] = { 5'd14,	5'd8,	5'd6,	5'd12};
		rom[ 1330 ] = { 5'd4,	5'd8,	5'd6,	5'd12};
		rom[ 1331 ] = { 5'd16,	5'd5,	5'd5,	5'd15};
		rom[ 1332 ] = { 5'd3,	5'd5,	5'd5,	5'd15};
		rom[ 1333 ] = { 5'd18,	5'd4,	5'd6,	5'd9};
		rom[ 1334 ] = { 5'd1,	5'd7,	5'd6,	5'd15};
		rom[ 1335 ] = { 5'd11,	5'd15,	5'd12,	5'd8};
		rom[ 1336 ] = { 5'd0,	5'd2,	5'd24,	5'd4};
		rom[ 1337 ] = { 5'd15,	5'd1,	5'd2,	5'd19};
		rom[ 1338 ] = { 5'd7,	5'd1,	5'd2,	5'd19};
		rom[ 1339 ] = { 5'd22,	5'd1,	5'd2,	5'd20};
		rom[ 1340 ] = { 5'd0,	5'd1,	5'd2,	5'd20};
		rom[ 1341 ] = { 5'd18,	5'd11,	5'd6,	5'd12};
		rom[ 1342 ] = { 5'd0,	5'd11,	5'd6,	5'd12};
		rom[ 1343 ] = { 5'd3,	5'd6,	5'd18,	5'd14};
		rom[ 1344 ] = { 5'd6,	5'd10,	5'd7,	5'd8};
		rom[ 1345 ] = { 5'd7,	5'd9,	5'd12,	5'd12};
		rom[ 1346 ] = { 5'd2,	5'd18,	5'd18,	5'd5};
		rom[ 1347 ] = { 5'd4,	5'd21,	5'd20,	5'd3};
		rom[ 1348 ] = { 5'd9,	5'd12,	5'd6,	5'd12};
		rom[ 1349 ] = { 5'd4,	5'd6,	5'd18,	5'd3};
		rom[ 1350 ] = { 5'd3,	5'd6,	5'd18,	5'd3};
		rom[ 1351 ] = { 5'd18,	5'd4,	5'd6,	5'd9};
		rom[ 1352 ] = { 5'd2,	5'd12,	5'd9,	5'd6};
		rom[ 1353 ] = { 5'd4,	5'd14,	5'd18,	5'd4};
		rom[ 1354 ] = { 5'd7,	5'd7,	5'd6,	5'd14};
		rom[ 1355 ] = { 5'd7,	5'd13,	5'd12,	5'd6};
		rom[ 1356 ] = { 5'd6,	5'd7,	5'd12,	5'd9};
		rom[ 1357 ] = { 5'd12,	5'd12,	5'd6,	5'd6};
		rom[ 1358 ] = { 5'd0,	5'd2,	5'd4,	5'd10};
		rom[ 1359 ] = { 5'd8,	5'd0,	5'd9,	5'd6};
		rom[ 1360 ] = { 5'd2,	5'd9,	5'd12,	5'd6};
		rom[ 1361 ] = { 5'd13,	5'd10,	5'd6,	5'd9};
		rom[ 1362 ] = { 5'd5,	5'd10,	5'd6,	5'd9};
		rom[ 1363 ] = { 5'd9,	5'd15,	5'd9,	5'd6};
		rom[ 1364 ] = { 5'd5,	5'd16,	5'd12,	5'd6};
		rom[ 1365 ] = { 5'd3,	5'd2,	5'd20,	5'd3};
		rom[ 1366 ] = { 5'd2,	5'd5,	5'd12,	5'd6};
		rom[ 1367 ] = { 5'd11,	5'd0,	5'd3,	5'd24};
		rom[ 1368 ] = { 5'd3,	5'd16,	5'd15,	5'd4};
		rom[ 1369 ] = { 5'd9,	5'd12,	5'd6,	5'd12};
		rom[ 1370 ] = { 5'd1,	5'd15,	5'd12,	5'd8};
		rom[ 1371 ] = { 5'd15,	5'd10,	5'd8,	5'd14};
		rom[ 1372 ] = { 5'd1,	5'd9,	5'd8,	5'd14};
		rom[ 1373 ] = { 5'd9,	5'd11,	5'd9,	5'd10};
		rom[ 1374 ] = { 5'd6,	5'd7,	5'd12,	5'd6};
		rom[ 1375 ] = { 5'd10,	5'd15,	5'd6,	5'd9};
		rom[ 1376 ] = { 5'd7,	5'd8,	5'd9,	5'd7};
		rom[ 1377 ] = { 5'd10,	5'd4,	5'd8,	5'd10};
		rom[ 1378 ] = { 5'd4,	5'd6,	5'd6,	5'd9};
		rom[ 1379 ] = { 5'd0,	5'd6,	5'd24,	5'd12};
		rom[ 1380 ] = { 5'd3,	5'd7,	5'd6,	5'd14};
		rom[ 1381 ] = { 5'd19,	5'd8,	5'd5,	5'd8};
		rom[ 1382 ] = { 5'd0,	5'd8,	5'd5,	5'd8};
		rom[ 1383 ] = { 5'd17,	5'd3,	5'd6,	5'd6};
		rom[ 1384 ] = { 5'd1,	5'd3,	5'd6,	5'd6};
		rom[ 1385 ] = { 5'd18,	5'd2,	5'd6,	5'd9};
		rom[ 1386 ] = { 5'd0,	5'd2,	5'd6,	5'd9};
		rom[ 1387 ] = { 5'd3,	5'd3,	5'd18,	5'd6};
		rom[ 1388 ] = { 5'd2,	5'd3,	5'd9,	5'd6};
		rom[ 1389 ] = { 5'd9,	5'd3,	5'd10,	5'd8};
		rom[ 1390 ] = { 5'd5,	5'd3,	5'd10,	5'd8};
		rom[ 1391 ] = { 5'd10,	5'd11,	5'd6,	5'd12};
		rom[ 1392 ] = { 5'd8,	5'd11,	5'd6,	5'd11};
		rom[ 1393 ] = { 5'd7,	5'd8,	5'd10,	5'd4};
		rom[ 1394 ] = { 5'd9,	5'd6,	5'd6,	5'd7};
		rom[ 1395 ] = { 5'd5,	5'd18,	5'd18,	5'd3};
		rom[ 1396 ] = { 5'd8,	5'd4,	5'd6,	5'd9};
		rom[ 1397 ] = { 5'd8,	5'd1,	5'd9,	5'd7};
		rom[ 1398 ] = { 5'd6,	5'd11,	5'd6,	5'd6};
		rom[ 1399 ] = { 5'd14,	5'd12,	5'd4,	5'd11};
		rom[ 1400 ] = { 5'd6,	5'd12,	5'd4,	5'd11};
		rom[ 1401 ] = { 5'd8,	5'd0,	5'd12,	5'd18};
		rom[ 1402 ] = { 5'd2,	5'd12,	5'd10,	5'd5};
		rom[ 1403 ] = { 5'd2,	5'd20,	5'd22,	5'd3};
		rom[ 1404 ] = { 5'd0,	5'd4,	5'd2,	5'd20};
		rom[ 1405 ] = { 5'd0,	5'd2,	5'd24,	5'd4};
		rom[ 1406 ] = { 5'd7,	5'd8,	5'd10,	5'd4};
		rom[ 1407 ] = { 5'd6,	5'd7,	5'd8,	5'd10};
		rom[ 1408 ] = { 5'd14,	5'd0,	5'd6,	5'd14};
		rom[ 1409 ] = { 5'd4,	5'd11,	5'd5,	5'd8};
		rom[ 1410 ] = { 5'd2,	5'd0,	5'd20,	5'd9};
		rom[ 1411 ] = { 5'd6,	5'd7,	5'd12,	5'd8};
		rom[ 1412 ] = { 5'd9,	5'd17,	5'd6,	5'd6};
		rom[ 1413 ] = { 5'd7,	5'd10,	5'd10,	5'd4};
		rom[ 1414 ] = { 5'd6,	5'd5,	5'd12,	5'd9};
		rom[ 1415 ] = { 5'd5,	5'd11,	5'd6,	5'd8};
		rom[ 1416 ] = { 5'd18,	5'd4,	5'd4,	5'd17};
		rom[ 1417 ] = { 5'd0,	5'd0,	5'd6,	5'd6};
		rom[ 1418 ] = { 5'd18,	5'd4,	5'd4,	5'd17};
		rom[ 1419 ] = { 5'd2,	5'd4,	5'd4,	5'd17};
		rom[ 1420 ] = { 5'd5,	5'd18,	5'd19,	5'd3};
		rom[ 1421 ] = { 5'd11,	5'd0,	5'd2,	5'd18};
		rom[ 1422 ] = { 5'd15,	5'd4,	5'd2,	5'd18};
		rom[ 1423 ] = { 5'd7,	5'd4,	5'd2,	5'd18};
		rom[ 1424 ] = { 5'd7,	5'd11,	5'd10,	5'd8};
		rom[ 1425 ] = { 5'd10,	5'd6,	5'd4,	5'd9};
		rom[ 1426 ] = { 5'd10,	5'd0,	5'd6,	5'd9};
		rom[ 1427 ] = { 5'd2,	5'd9,	5'd16,	5'd8};
		rom[ 1428 ] = { 5'd14,	5'd15,	5'd6,	5'd9};
		rom[ 1429 ] = { 5'd8,	5'd7,	5'd6,	5'd9};
		rom[ 1430 ] = { 5'd14,	5'd15,	5'd6,	5'd9};
		rom[ 1431 ] = { 5'd3,	5'd12,	5'd12,	5'd6};
		rom[ 1432 ] = { 5'd14,	5'd12,	5'd9,	5'd6};
		rom[ 1433 ] = { 5'd1,	5'd12,	5'd9,	5'd6};
		rom[ 1434 ] = { 5'd3,	5'd7,	5'd18,	5'd3};
		rom[ 1435 ] = { 5'd1,	5'd7,	5'd22,	5'd6};
		rom[ 1436 ] = { 5'd18,	5'd4,	5'd6,	5'd6};
		rom[ 1437 ] = { 5'd0,	5'd4,	5'd6,	5'd6};
		rom[ 1438 ] = { 5'd5,	5'd11,	5'd16,	5'd6};
		rom[ 1439 ] = { 5'd6,	5'd16,	5'd9,	5'd4};
		rom[ 1440 ] = { 5'd14,	5'd15,	5'd6,	5'd9};
		rom[ 1441 ] = { 5'd4,	5'd15,	5'd6,	5'd9};
		rom[ 1442 ] = { 5'd15,	5'd1,	5'd6,	5'd23};
		rom[ 1443 ] = { 5'd0,	5'd21,	5'd24,	5'd3};
		rom[ 1444 ] = { 5'd0,	5'd20,	5'd24,	5'd4};
		rom[ 1445 ] = { 5'd3,	5'd1,	5'd6,	5'd23};
		rom[ 1446 ] = { 5'd3,	5'd17,	5'd18,	5'd3};
		rom[ 1447 ] = { 5'd0,	5'd16,	5'd18,	5'd3};
		rom[ 1448 ] = { 5'd1,	5'd16,	5'd22,	5'd4};
		rom[ 1449 ] = { 5'd0,	5'd16,	5'd9,	5'd6};
		rom[ 1450 ] = { 5'd2,	5'd10,	5'd21,	5'd3};
		rom[ 1451 ] = { 5'd2,	5'd18,	5'd12,	5'd6};
		rom[ 1452 ] = { 5'd0,	5'd5,	5'd24,	5'd4};
		rom[ 1453 ] = { 5'd10,	5'd2,	5'd4,	5'd15};
		rom[ 1454 ] = { 5'd10,	5'd7,	5'd6,	5'd12};
		rom[ 1455 ] = { 5'd6,	5'd6,	5'd6,	5'd9};
		rom[ 1456 ] = { 5'd11,	5'd0,	5'd6,	5'd9};
		rom[ 1457 ] = { 5'd9,	5'd7,	5'd6,	5'd9};
		rom[ 1458 ] = { 5'd2,	5'd1,	5'd20,	5'd3};
		rom[ 1459 ] = { 5'd1,	5'd18,	5'd12,	5'd6};
		rom[ 1460 ] = { 5'd13,	5'd2,	5'd4,	5'd13};
		rom[ 1461 ] = { 5'd6,	5'd7,	5'd12,	5'd4};
		rom[ 1462 ] = { 5'd10,	5'd1,	5'd4,	5'd13};
		rom[ 1463 ] = { 5'd6,	5'd0,	5'd3,	5'd18};
		rom[ 1464 ] = { 5'd14,	5'd3,	5'd10,	5'd5};
		rom[ 1465 ] = { 5'd6,	5'd15,	5'd12,	5'd8};
		rom[ 1466 ] = { 5'd9,	5'd10,	5'd6,	5'd9};
		rom[ 1467 ] = { 5'd8,	5'd3,	5'd4,	5'd9};
		rom[ 1468 ] = { 5'd17,	5'd0,	5'd6,	5'd14};
		rom[ 1469 ] = { 5'd1,	5'd0,	5'd6,	5'd14};
		rom[ 1470 ] = { 5'd14,	5'd0,	5'd6,	5'd16};
		rom[ 1471 ] = { 5'd7,	5'd4,	5'd4,	5'd10};
		rom[ 1472 ] = { 5'd3,	5'd17,	5'd18,	5'd6};
		rom[ 1473 ] = { 5'd1,	5'd20,	5'd22,	5'd4};
		rom[ 1474 ] = { 5'd14,	5'd3,	5'd10,	5'd5};
		rom[ 1475 ] = { 5'd0,	5'd3,	5'd10,	5'd5};
		rom[ 1476 ] = { 5'd12,	5'd6,	5'd12,	5'd16};
		rom[ 1477 ] = { 5'd0,	5'd6,	5'd12,	5'd16};
		rom[ 1478 ] = { 5'd10,	5'd9,	5'd5,	5'd15};
		rom[ 1479 ] = { 5'd1,	5'd18,	5'd21,	5'd2};
		rom[ 1480 ] = { 5'd15,	5'd0,	5'd9,	5'd6};
		rom[ 1481 ] = { 5'd6,	5'd1,	5'd12,	5'd4};
		rom[ 1482 ] = { 5'd6,	5'd0,	5'd12,	5'd12};
		rom[ 1483 ] = { 5'd8,	5'd10,	5'd8,	5'd12};
		rom[ 1484 ] = { 5'd14,	5'd16,	5'd10,	5'd8};
		rom[ 1485 ] = { 5'd0,	5'd16,	5'd10,	5'd8};
		rom[ 1486 ] = { 5'd10,	5'd12,	5'd12,	5'd5};
		rom[ 1487 ] = { 5'd6,	5'd16,	5'd10,	5'd8};
		rom[ 1488 ] = { 5'd7,	5'd6,	5'd12,	5'd6};
		rom[ 1489 ] = { 5'd9,	5'd6,	5'd4,	5'd18};
		rom[ 1490 ] = { 5'd10,	5'd9,	5'd6,	5'd14};
		rom[ 1491 ] = { 5'd8,	5'd9,	5'd6,	5'd14};
		rom[ 1492 ] = { 5'd7,	5'd4,	5'd11,	5'd12};
		rom[ 1493 ] = { 5'd4,	5'd8,	5'd6,	5'd16};
		rom[ 1494 ] = { 5'd17,	5'd3,	5'd4,	5'd21};
		rom[ 1495 ] = { 5'd3,	5'd3,	5'd4,	5'd21};
		rom[ 1496 ] = { 5'd10,	5'd1,	5'd8,	5'd18};
		rom[ 1497 ] = { 5'd2,	5'd5,	5'd16,	5'd8};
		rom[ 1498 ] = { 5'd3,	5'd6,	5'd18,	5'd12};
		rom[ 1499 ] = { 5'd4,	5'd10,	5'd16,	5'd12};
		rom[ 1500 ] = { 5'd15,	5'd4,	5'd8,	5'd20};
		rom[ 1501 ] = { 5'd7,	5'd2,	5'd9,	5'd6};
		rom[ 1502 ] = { 5'd15,	5'd4,	5'd8,	5'd20};
		rom[ 1503 ] = { 5'd1,	5'd4,	5'd8,	5'd20};
		rom[ 1504 ] = { 5'd11,	5'd8,	5'd8,	5'd14};
		rom[ 1505 ] = { 5'd5,	5'd8,	5'd8,	5'd14};
		rom[ 1506 ] = { 5'd10,	5'd13,	5'd5,	5'd8};
		rom[ 1507 ] = { 5'd4,	5'd13,	5'd7,	5'd9};
		rom[ 1508 ] = { 5'd0,	5'd13,	5'd24,	5'd10};
		rom[ 1509 ] = { 5'd4,	5'd2,	5'd8,	5'd11};
		rom[ 1510 ] = { 5'd10,	5'd2,	5'd8,	5'd16};
		rom[ 1511 ] = { 5'd0,	5'd2,	5'd24,	5'd6};
		rom[ 1512 ] = { 5'd6,	5'd0,	5'd12,	5'd9};
		rom[ 1513 ] = { 5'd1,	5'd2,	5'd12,	5'd12};
		rom[ 1514 ] = { 5'd18,	5'd5,	5'd6,	5'd9};
		rom[ 1515 ] = { 5'd4,	5'd3,	5'd8,	5'd10};
		rom[ 1516 ] = { 5'd6,	5'd21,	5'd18,	5'd3};
		rom[ 1517 ] = { 5'd1,	5'd10,	5'd18,	5'd2};
		rom[ 1518 ] = { 5'd1,	5'd10,	5'd22,	5'd3};
		rom[ 1519 ] = { 5'd2,	5'd8,	5'd12,	5'd9};
		rom[ 1520 ] = { 5'd12,	5'd8,	5'd12,	5'd6};
		rom[ 1521 ] = { 5'd0,	5'd8,	5'd12,	5'd6};
		rom[ 1522 ] = { 5'd10,	5'd15,	5'd6,	5'd9};
		rom[ 1523 ] = { 5'd7,	5'd13,	5'd9,	5'd6};
		rom[ 1524 ] = { 5'd9,	5'd8,	5'd7,	5'd12};
		rom[ 1525 ] = { 5'd4,	5'd13,	5'd9,	5'd6};
		rom[ 1526 ] = { 5'd6,	5'd15,	5'd18,	5'd4};
		rom[ 1527 ] = { 5'd5,	5'd4,	5'd4,	5'd16};
		rom[ 1528 ] = { 5'd10,	5'd15,	5'd6,	5'd9};
		rom[ 1529 ] = { 5'd8,	5'd15,	5'd6,	5'd9};
		rom[ 1530 ] = { 5'd9,	5'd11,	5'd12,	5'd10};
		rom[ 1531 ] = { 5'd3,	5'd6,	5'd14,	5'd6};
		rom[ 1532 ] = { 5'd4,	5'd2,	5'd17,	5'd8};
		rom[ 1533 ] = { 5'd6,	5'd2,	5'd12,	5'd21};
		rom[ 1534 ] = { 5'd8,	5'd1,	5'd9,	5'd9};
		rom[ 1535 ] = { 5'd0,	5'd7,	5'd24,	5'd3};
		rom[ 1536 ] = { 5'd11,	5'd6,	5'd9,	5'd10};
		rom[ 1537 ] = { 5'd2,	5'd11,	5'd18,	5'd3};
		rom[ 1538 ] = { 5'd8,	5'd16,	5'd9,	5'd4};
		rom[ 1539 ] = { 5'd0,	5'd0,	5'd9,	5'd6};
		rom[ 1540 ] = { 5'd0,	5'd11,	5'd24,	5'd6};
		rom[ 1541 ] = { 5'd2,	5'd9,	5'd20,	5'd6};
		rom[ 1542 ] = { 5'd4,	5'd5,	5'd16,	5'd12};
		rom[ 1543 ] = { 5'd10,	5'd2,	5'd4,	5'd15};
		rom[ 1544 ] = { 5'd7,	5'd3,	5'd10,	5'd4};
		rom[ 1545 ] = { 5'd9,	5'd15,	5'd6,	5'd8};
		rom[ 1546 ] = { 5'd17,	5'd0,	5'd7,	5'd10};
		rom[ 1547 ] = { 5'd0,	5'd0,	5'd7,	5'd10};
		rom[ 1548 ] = { 5'd16,	5'd1,	5'd6,	5'd12};
		rom[ 1549 ] = { 5'd1,	5'd0,	5'd19,	5'd8};
		rom[ 1550 ] = { 5'd12,	5'd2,	5'd9,	5'd4};
		rom[ 1551 ] = { 5'd3,	5'd2,	5'd9,	5'd4};
		rom[ 1552 ] = { 5'd12,	5'd2,	5'd10,	5'd6};
		rom[ 1553 ] = { 5'd3,	5'd4,	5'd18,	5'd2};
		rom[ 1554 ] = { 5'd12,	5'd1,	5'd4,	5'd9};
		rom[ 1555 ] = { 5'd8,	5'd1,	5'd4,	5'd9};
		rom[ 1556 ] = { 5'd10,	5'd5,	5'd8,	5'd10};
		rom[ 1557 ] = { 5'd6,	5'd4,	5'd12,	5'd13};
		rom[ 1558 ] = { 5'd13,	5'd5,	5'd6,	5'd6};
		rom[ 1559 ] = { 5'd1,	5'd5,	5'd12,	5'd3};
		rom[ 1560 ] = { 5'd7,	5'd5,	5'd10,	5'd6};
		rom[ 1561 ] = { 5'd2,	5'd0,	5'd21,	5'd5};
		rom[ 1562 ] = { 5'd0,	5'd8,	5'd9,	5'd9};
		rom[ 1563 ] = { 5'd9,	5'd6,	5'd6,	5'd9};
		rom[ 1564 ] = { 5'd0,	5'd3,	5'd6,	5'd7};
		rom[ 1565 ] = { 5'd9,	5'd18,	5'd12,	5'd6};
		rom[ 1566 ] = { 5'd2,	5'd8,	5'd20,	5'd6};
		rom[ 1567 ] = { 5'd13,	5'd2,	5'd10,	5'd4};
		rom[ 1568 ] = { 5'd4,	5'd5,	5'd5,	5'd18};
		rom[ 1569 ] = { 5'd20,	5'd4,	5'd4,	5'd9};
		rom[ 1570 ] = { 5'd8,	5'd6,	5'd8,	5'd14};
		rom[ 1571 ] = { 5'd0,	5'd1,	5'd24,	5'd6};
		rom[ 1572 ] = { 5'd0,	5'd4,	5'd4,	5'd9};
		rom[ 1573 ] = { 5'd3,	5'd6,	5'd18,	5'd3};
		rom[ 1574 ] = { 5'd3,	5'd17,	5'd16,	5'd6};
		rom[ 1575 ] = { 5'd13,	5'd6,	5'd6,	5'd9};
		rom[ 1576 ] = { 5'd5,	5'd6,	5'd14,	5'd6};
		rom[ 1577 ] = { 5'd13,	5'd5,	5'd8,	5'd10};
		rom[ 1578 ] = { 5'd2,	5'd2,	5'd20,	5'd3};
		rom[ 1579 ] = { 5'd9,	5'd2,	5'd9,	5'd6};
		rom[ 1580 ] = { 5'd8,	5'd6,	5'd6,	5'd9};
		rom[ 1581 ] = { 5'd12,	5'd3,	5'd4,	5'd11};
		rom[ 1582 ] = { 5'd8,	5'd3,	5'd4,	5'd11};
		rom[ 1583 ] = { 5'd8,	5'd3,	5'd8,	5'd10};
		rom[ 1584 ] = { 5'd11,	5'd1,	5'd2,	5'd18};
		rom[ 1585 ] = { 5'd9,	5'd2,	5'd9,	5'd6};
		rom[ 1586 ] = { 5'd0,	5'd2,	5'd19,	5'd3};
		rom[ 1587 ] = { 5'd9,	5'd14,	5'd9,	5'd6};
		rom[ 1588 ] = { 5'd1,	5'd8,	5'd18,	5'd5};
		rom[ 1589 ] = { 5'd12,	5'd0,	5'd6,	5'd9};
		rom[ 1590 ] = { 5'd6,	5'd0,	5'd6,	5'd9};
		rom[ 1591 ] = { 5'd13,	5'd6,	5'd4,	5'd15};
		rom[ 1592 ] = { 5'd1,	5'd5,	5'd18,	5'd3};
		rom[ 1593 ] = { 5'd9,	5'd7,	5'd14,	5'd6};
		rom[ 1594 ] = { 5'd2,	5'd16,	5'd18,	5'd3};
		rom[ 1595 ] = { 5'd15,	5'd17,	5'd9,	5'd6};
		rom[ 1596 ] = { 5'd0,	5'd8,	5'd12,	5'd6};
		rom[ 1597 ] = { 5'd9,	5'd13,	5'd7,	5'd8};
		rom[ 1598 ] = { 5'd2,	5'd17,	5'd20,	5'd3};
		rom[ 1599 ] = { 5'd15,	5'd17,	5'd9,	5'd6};
		rom[ 1600 ] = { 5'd4,	5'd0,	5'd15,	5'd4};
		rom[ 1601 ] = { 5'd17,	5'd2,	5'd6,	5'd6};
		rom[ 1602 ] = { 5'd0,	5'd3,	5'd6,	5'd9};
		rom[ 1603 ] = { 5'd15,	5'd17,	5'd9,	5'd6};
		rom[ 1604 ] = { 5'd0,	5'd17,	5'd9,	5'd6};
		rom[ 1605 ] = { 5'd9,	5'd18,	5'd12,	5'd6};
		rom[ 1606 ] = { 5'd3,	5'd15,	5'd6,	5'd9};
		rom[ 1607 ] = { 5'd16,	5'd13,	5'd8,	5'd10};
		rom[ 1608 ] = { 5'd0,	5'd14,	5'd24,	5'd4};
		rom[ 1609 ] = { 5'd13,	5'd18,	5'd6,	5'd6};
		rom[ 1610 ] = { 5'd0,	5'd13,	5'd8,	5'd10};
		rom[ 1611 ] = { 5'd0,	5'd14,	5'd24,	5'd6};
		rom[ 1612 ] = { 5'd5,	5'd2,	5'd12,	5'd8};
		rom[ 1613 ] = { 5'd8,	5'd9,	5'd9,	5'd6};
		rom[ 1614 ] = { 5'd4,	5'd3,	5'd16,	5'd4};
		rom[ 1615 ] = { 5'd10,	5'd2,	5'd4,	5'd10};
		rom[ 1616 ] = { 5'd8,	5'd4,	5'd5,	5'd8};
		rom[ 1617 ] = { 5'd11,	5'd5,	5'd9,	5'd12};
		rom[ 1618 ] = { 5'd4,	5'd5,	5'd9,	5'd12};
		rom[ 1619 ] = { 5'd14,	5'd6,	5'd6,	5'd9};
		rom[ 1620 ] = { 5'd2,	5'd4,	5'd20,	5'd12};
		rom[ 1621 ] = { 5'd4,	5'd4,	5'd17,	5'd16};
		rom[ 1622 ] = { 5'd8,	5'd7,	5'd7,	5'd6};
		rom[ 1623 ] = { 5'd1,	5'd9,	5'd23,	5'd2};
		rom[ 1624 ] = { 5'd7,	5'd0,	5'd6,	5'd9};
		rom[ 1625 ] = { 5'd13,	5'd3,	5'd4,	5'd9};
		rom[ 1626 ] = { 5'd8,	5'd1,	5'd6,	5'd13};
		rom[ 1627 ] = { 5'd4,	5'd22,	5'd18,	5'd2};
		rom[ 1628 ] = { 5'd3,	5'd10,	5'd9,	5'd6};
		rom[ 1629 ] = { 5'd14,	5'd0,	5'd2,	5'd24};
		rom[ 1630 ] = { 5'd8,	5'd0,	5'd2,	5'd24};
		rom[ 1631 ] = { 5'd3,	5'd2,	5'd18,	5'd10};
		rom[ 1632 ] = { 5'd4,	5'd13,	5'd15,	5'd6};
		rom[ 1633 ] = { 5'd3,	5'd21,	5'd18,	5'd3};
		rom[ 1634 ] = { 5'd9,	5'd1,	5'd4,	5'd11};
		rom[ 1635 ] = { 5'd9,	5'd7,	5'd10,	5'd4};
		rom[ 1636 ] = { 5'd7,	5'd0,	5'd10,	5'd18};
		rom[ 1637 ] = { 5'd12,	5'd1,	5'd6,	5'd16};
		rom[ 1638 ] = { 5'd6,	5'd1,	5'd6,	5'd16};
		rom[ 1639 ] = { 5'd18,	5'd2,	5'd6,	5'd6};
		rom[ 1640 ] = { 5'd3,	5'd5,	5'd18,	5'd2};
		rom[ 1641 ] = { 5'd18,	5'd2,	5'd6,	5'd6};
		rom[ 1642 ] = { 5'd0,	5'd2,	5'd6,	5'd6};
		rom[ 1643 ] = { 5'd13,	5'd11,	5'd11,	5'd6};
		rom[ 1644 ] = { 5'd5,	5'd7,	5'd10,	5'd4};
		rom[ 1645 ] = { 5'd11,	5'd9,	5'd10,	5'd7};
		rom[ 1646 ] = { 5'd3,	5'd9,	5'd10,	5'd7};
		rom[ 1647 ] = { 5'd16,	5'd4,	5'd6,	5'd6};
		rom[ 1648 ] = { 5'd5,	5'd6,	5'd10,	5'd8};
		rom[ 1649 ] = { 5'd7,	5'd21,	5'd16,	5'd3};
		rom[ 1650 ] = { 5'd1,	5'd21,	5'd16,	5'd3};
		rom[ 1651 ] = { 5'd2,	5'd5,	5'd22,	5'd14};
		rom[ 1652 ] = { 5'd3,	5'd10,	5'd8,	5'd10};
		rom[ 1653 ] = { 5'd17,	5'd0,	5'd6,	5'd12};
		rom[ 1654 ] = { 5'd5,	5'd2,	5'd6,	5'd18};
		rom[ 1655 ] = { 5'd13,	5'd0,	5'd6,	5'd9};
		rom[ 1656 ] = { 5'd0,	5'd12,	5'd7,	5'd9};
		rom[ 1657 ] = { 5'd15,	5'd13,	5'd8,	5'd10};
		rom[ 1658 ] = { 5'd1,	5'd0,	5'd6,	5'd12};
		rom[ 1659 ] = { 5'd12,	5'd1,	5'd3,	5'd12};
		rom[ 1660 ] = { 5'd1,	5'd13,	5'd8,	5'd10};
		rom[ 1661 ] = { 5'd3,	5'd21,	5'd19,	5'd2};
		rom[ 1662 ] = { 5'd6,	5'd3,	5'd4,	5'd13};
		rom[ 1663 ] = { 5'd5,	5'd10,	5'd18,	5'd3};
		rom[ 1664 ] = { 5'd9,	5'd3,	5'd5,	5'd12};
		rom[ 1665 ] = { 5'd11,	5'd2,	5'd4,	5'd15};
		rom[ 1666 ] = { 5'd4,	5'd1,	5'd16,	5'd4};
		rom[ 1667 ] = { 5'd6,	5'd0,	5'd18,	5'd3};
		rom[ 1668 ] = { 5'd5,	5'd1,	5'd10,	5'd8};
		rom[ 1669 ] = { 5'd11,	5'd18,	5'd12,	5'd6};
		rom[ 1670 ] = { 5'd5,	5'd15,	5'd12,	5'd3};
		rom[ 1671 ] = { 5'd1,	5'd10,	5'd22,	5'd4};
		rom[ 1672 ] = { 5'd7,	5'd9,	5'd9,	5'd6};
		rom[ 1673 ] = { 5'd6,	5'd11,	5'd12,	5'd5};
		rom[ 1674 ] = { 5'd6,	5'd7,	5'd10,	5'd7};
		rom[ 1675 ] = { 5'd11,	5'd2,	5'd8,	5'd10};
		rom[ 1676 ] = { 5'd5,	5'd2,	5'd8,	5'd10};
		rom[ 1677 ] = { 5'd6,	5'd4,	5'd18,	5'd6};
		rom[ 1678 ] = { 5'd0,	5'd5,	5'd10,	5'd9};
		rom[ 1679 ] = { 5'd2,	5'd7,	5'd21,	5'd6};
		rom[ 1680 ] = { 5'd0,	5'd4,	5'd22,	5'd16};
		rom[ 1681 ] = { 5'd9,	5'd0,	5'd6,	5'd22};
		rom[ 1682 ] = { 5'd9,	5'd1,	5'd3,	5'd12};
		rom[ 1683 ] = { 5'd12,	5'd0,	5'd12,	5'd18};
		rom[ 1684 ] = { 5'd0,	5'd0,	5'd12,	5'd18};
		rom[ 1685 ] = { 5'd1,	5'd1,	5'd22,	5'd4};
		rom[ 1686 ] = { 5'd3,	5'd0,	5'd18,	5'd4};
		rom[ 1687 ] = { 5'd2,	5'd5,	5'd22,	5'd6};
		rom[ 1688 ] = { 5'd5,	5'd0,	5'd6,	5'd9};
		rom[ 1689 ] = { 5'd10,	5'd14,	5'd6,	5'd9};
		rom[ 1690 ] = { 5'd8,	5'd14,	5'd6,	5'd9};
		rom[ 1691 ] = { 5'd5,	5'd18,	5'd18,	5'd3};
		rom[ 1692 ] = { 5'd6,	5'd0,	5'd6,	5'd13};
		rom[ 1693 ] = { 5'd7,	5'd4,	5'd12,	5'd4};
		rom[ 1694 ] = { 5'd5,	5'd2,	5'd12,	5'd6};
		rom[ 1695 ] = { 5'd4,	5'd1,	5'd18,	5'd3};
		rom[ 1696 ] = { 5'd0,	5'd8,	5'd6,	5'd12};
		rom[ 1697 ] = { 5'd9,	5'd15,	5'd6,	5'd9};
		rom[ 1698 ] = { 5'd9,	5'd10,	5'd6,	5'd13};
		rom[ 1699 ] = { 5'd6,	5'd17,	5'd18,	5'd2};
		rom[ 1700 ] = { 5'd9,	5'd4,	5'd6,	5'd9};
		rom[ 1701 ] = { 5'd10,	5'd0,	5'd6,	5'd9};
		rom[ 1702 ] = { 5'd5,	5'd6,	5'd10,	5'd8};
		rom[ 1703 ] = { 5'd14,	5'd9,	5'd5,	5'd8};
		rom[ 1704 ] = { 5'd5,	5'd9,	5'd5,	5'd8};
		rom[ 1705 ] = { 5'd14,	5'd11,	5'd9,	5'd6};
		rom[ 1706 ] = { 5'd0,	5'd2,	5'd23,	5'd15};
		rom[ 1707 ] = { 5'd16,	5'd0,	5'd8,	5'd12};
		rom[ 1708 ] = { 5'd4,	5'd15,	5'd6,	5'd9};
		rom[ 1709 ] = { 5'd8,	5'd18,	5'd9,	5'd4};
		rom[ 1710 ] = { 5'd0,	5'd17,	5'd18,	5'd3};
		rom[ 1711 ] = { 5'd13,	5'd11,	5'd11,	5'd6};
		rom[ 1712 ] = { 5'd0,	5'd11,	5'd11,	5'd6};
		rom[ 1713 ] = { 5'd0,	5'd9,	5'd24,	5'd6};
		rom[ 1714 ] = { 5'd6,	5'd16,	5'd8,	5'd8};
		rom[ 1715 ] = { 5'd10,	5'd16,	5'd14,	5'd6};
		rom[ 1716 ] = { 5'd1,	5'd1,	5'd21,	5'd3};
		rom[ 1717 ] = { 5'd0,	5'd2,	5'd24,	5'd3};
		rom[ 1718 ] = { 5'd2,	5'd15,	5'd8,	5'd5};
		rom[ 1719 ] = { 5'd2,	5'd11,	5'd21,	5'd3};
		rom[ 1720 ] = { 5'd1,	5'd18,	5'd12,	5'd6};
		rom[ 1721 ] = { 5'd10,	5'd14,	5'd4,	5'd10};
		rom[ 1722 ] = { 5'd7,	5'd7,	5'd4,	5'd10};
		rom[ 1723 ] = { 5'd9,	5'd8,	5'd6,	5'd12};
		rom[ 1724 ] = { 5'd7,	5'd1,	5'd9,	5'd6};
		rom[ 1725 ] = { 5'd3,	5'd14,	5'd19,	5'd2};
		rom[ 1726 ] = { 5'd7,	5'd7,	5'd10,	5'd10};
		rom[ 1727 ] = { 5'd3,	5'd12,	5'd18,	5'd12};
		rom[ 1728 ] = { 5'd8,	5'd0,	5'd6,	5'd12};
		rom[ 1729 ] = { 5'd3,	5'd0,	5'd17,	5'd9};
		rom[ 1730 ] = { 5'd6,	5'd0,	5'd12,	5'd11};
		rom[ 1731 ] = { 5'd1,	5'd0,	5'd6,	5'd13};
		rom[ 1732 ] = { 5'd5,	5'd8,	5'd16,	5'd6};
		rom[ 1733 ] = { 5'd8,	5'd8,	5'd5,	5'd12};
		rom[ 1734 ] = { 5'd3,	5'd21,	5'd18,	5'd3};
		rom[ 1735 ] = { 5'd0,	5'd0,	5'd6,	5'd6};
		rom[ 1736 ] = { 5'd2,	5'd0,	5'd20,	5'd3};
		rom[ 1737 ] = { 5'd4,	5'd6,	5'd15,	5'd10};
		rom[ 1738 ] = { 5'd9,	5'd6,	5'd6,	5'd9};
		rom[ 1739 ] = { 5'd9,	5'd0,	5'd6,	5'd9};
		rom[ 1740 ] = { 5'd14,	5'd0,	5'd6,	5'd9};
		rom[ 1741 ] = { 5'd7,	5'd16,	5'd9,	5'd6};
		rom[ 1742 ] = { 5'd14,	5'd0,	5'd6,	5'd9};
		rom[ 1743 ] = { 5'd4,	5'd0,	5'd6,	5'd9};
		rom[ 1744 ] = { 5'd17,	5'd1,	5'd6,	5'd16};
		rom[ 1745 ] = { 5'd1,	5'd1,	5'd6,	5'd16};
		rom[ 1746 ] = { 5'd14,	5'd13,	5'd6,	5'd9};
		rom[ 1747 ] = { 5'd0,	5'd0,	5'd6,	5'd9};
		rom[ 1748 ] = { 5'd9,	5'd5,	5'd6,	5'd6};
		rom[ 1749 ] = { 5'd3,	5'd10,	5'd9,	5'd6};
		rom[ 1750 ] = { 5'd14,	5'd7,	5'd3,	5'd16};
		rom[ 1751 ] = { 5'd4,	5'd10,	5'd14,	5'd12};
		rom[ 1752 ] = { 5'd7,	5'd6,	5'd12,	5'd6};
		rom[ 1753 ] = { 5'd7,	5'd2,	5'd4,	5'd20};
		rom[ 1754 ] = { 5'd14,	5'd13,	5'd6,	5'd9};
		rom[ 1755 ] = { 5'd10,	5'd6,	5'd4,	5'd9};
		rom[ 1756 ] = { 5'd14,	5'd13,	5'd6,	5'd9};
		rom[ 1757 ] = { 5'd5,	5'd20,	5'd14,	5'd4};
		rom[ 1758 ] = { 5'd4,	5'd4,	5'd16,	5'd12};
		rom[ 1759 ] = { 5'd9,	5'd6,	5'd6,	5'd9};
		rom[ 1760 ] = { 5'd3,	5'd0,	5'd21,	5'd4};
		rom[ 1761 ] = { 5'd4,	5'd13,	5'd6,	5'd9};
		rom[ 1762 ] = { 5'd16,	5'd16,	5'd5,	5'd8};
		rom[ 1763 ] = { 5'd4,	5'd0,	5'd16,	5'd16};
		rom[ 1764 ] = { 5'd6,	5'd6,	5'd14,	5'd6};
		rom[ 1765 ] = { 5'd10,	5'd5,	5'd4,	5'd15};
		rom[ 1766 ] = { 5'd9,	5'd15,	5'd12,	5'd8};
		rom[ 1767 ] = { 5'd6,	5'd7,	5'd12,	5'd4};
		rom[ 1768 ] = { 5'd5,	5'd6,	5'd14,	5'd6};
		rom[ 1769 ] = { 5'd3,	5'd6,	5'd18,	5'd10};
		rom[ 1770 ] = { 5'd6,	5'd0,	5'd18,	5'd21};
		rom[ 1771 ] = { 5'd0,	5'd0,	5'd24,	5'd21};
		rom[ 1772 ] = { 5'd6,	5'd18,	5'd18,	5'd3};
		rom[ 1773 ] = { 5'd0,	5'd15,	5'd9,	5'd6};
		rom[ 1774 ] = { 5'd4,	5'd3,	5'd19,	5'd2};
		rom[ 1775 ] = { 5'd0,	5'd3,	5'd24,	5'd2};
		rom[ 1776 ] = { 5'd15,	5'd14,	5'd9,	5'd4};
		rom[ 1777 ] = { 5'd0,	5'd14,	5'd9,	5'd4};
		rom[ 1778 ] = { 5'd6,	5'd15,	5'd18,	5'd2};
		rom[ 1779 ] = { 5'd3,	5'd17,	5'd18,	5'd3};
		rom[ 1780 ] = { 5'd12,	5'd0,	5'd3,	5'd23};
		rom[ 1781 ] = { 5'd6,	5'd0,	5'd8,	5'd6};
		rom[ 1782 ] = { 5'd6,	5'd16,	5'd18,	5'd3};
		rom[ 1783 ] = { 5'd9,	5'd0,	5'd3,	5'd23};
		rom[ 1784 ] = { 5'd10,	5'd7,	5'd4,	5'd10};
		rom[ 1785 ] = { 5'd7,	5'd8,	5'd10,	5'd12};
		rom[ 1786 ] = { 5'd14,	5'd9,	5'd6,	5'd14};
		rom[ 1787 ] = { 5'd2,	5'd0,	5'd10,	5'd9};
		rom[ 1788 ] = { 5'd11,	5'd1,	5'd5,	5'd12};
		rom[ 1789 ] = { 5'd1,	5'd4,	5'd12,	5'd10};
		rom[ 1790 ] = { 5'd15,	5'd1,	5'd9,	5'd4};
		rom[ 1791 ] = { 5'd1,	5'd2,	5'd8,	5'd10};
		rom[ 1792 ] = { 5'd10,	5'd1,	5'd5,	5'd12};
		rom[ 1793 ] = { 5'd4,	5'd0,	5'd14,	5'd24};
		rom[ 1794 ] = { 5'd7,	5'd17,	5'd10,	5'd4};
		rom[ 1795 ] = { 5'd10,	5'd14,	5'd4,	5'd10};
		rom[ 1796 ] = { 5'd13,	5'd15,	5'd6,	5'd9};
		rom[ 1797 ] = { 5'd3,	5'd21,	5'd18,	5'd3};
		rom[ 1798 ] = { 5'd13,	5'd15,	5'd6,	5'd9};
		rom[ 1799 ] = { 5'd5,	5'd15,	5'd6,	5'd9};
		rom[ 1800 ] = { 5'd10,	5'd6,	5'd4,	5'd18};
		rom[ 1801 ] = { 5'd7,	5'd3,	5'd6,	5'd11};
		rom[ 1802 ] = { 5'd15,	5'd1,	5'd9,	5'd4};
		rom[ 1803 ] = { 5'd5,	5'd4,	5'd14,	5'd8};
		rom[ 1804 ] = { 5'd8,	5'd1,	5'd15,	5'd9};
		rom[ 1805 ] = { 5'd7,	5'd2,	5'd8,	5'd10};
		rom[ 1806 ] = { 5'd12,	5'd2,	5'd6,	5'd12};
		rom[ 1807 ] = { 5'd6,	5'd2,	5'd6,	5'd12};
		rom[ 1808 ] = { 5'd7,	5'd7,	5'd12,	5'd4};
		rom[ 1809 ] = { 5'd6,	5'd3,	5'd12,	5'd10};
		rom[ 1810 ] = { 5'd5,	5'd6,	5'd16,	5'd6};
		rom[ 1811 ] = { 5'd3,	5'd1,	5'd18,	5'd9};
		rom[ 1812 ] = { 5'd3,	5'd8,	5'd18,	5'd5};
		rom[ 1813 ] = { 5'd0,	5'd0,	5'd24,	5'd22};
		rom[ 1814 ] = { 5'd14,	5'd16,	5'd9,	5'd6};
		rom[ 1815 ] = { 5'd0,	5'd16,	5'd24,	5'd8};
		rom[ 1816 ] = { 5'd1,	5'd19,	5'd22,	5'd4};
		rom[ 1817 ] = { 5'd1,	5'd16,	5'd9,	5'd6};
		rom[ 1818 ] = { 5'd7,	5'd8,	5'd10,	5'd4};
		rom[ 1819 ] = { 5'd9,	5'd15,	5'd6,	5'd9};
		rom[ 1820 ] = { 5'd10,	5'd18,	5'd12,	5'd6};
		rom[ 1821 ] = { 5'd2,	5'd18,	5'd12,	5'd6};
		rom[ 1822 ] = { 5'd8,	5'd3,	5'd16,	5'd9};
		rom[ 1823 ] = { 5'd0,	5'd5,	5'd10,	5'd6};
		rom[ 1824 ] = { 5'd5,	5'd5,	5'd18,	5'd3};
		rom[ 1825 ] = { 5'd2,	5'd6,	5'd9,	5'd6};
		rom[ 1826 ] = { 5'd14,	5'd2,	5'd10,	5'd9};
		rom[ 1827 ] = { 5'd3,	5'd6,	5'd18,	5'd3};
		rom[ 1828 ] = { 5'd9,	5'd2,	5'd15,	5'd6};
		rom[ 1829 ] = { 5'd4,	5'd8,	5'd15,	5'd6};
		rom[ 1830 ] = { 5'd0,	5'd5,	5'd24,	5'd4};
		rom[ 1831 ] = { 5'd7,	5'd8,	5'd6,	5'd12};
		rom[ 1832 ] = { 5'd11,	5'd0,	5'd6,	5'd9};
		rom[ 1833 ] = { 5'd0,	5'd12,	5'd6,	5'd12};
		rom[ 1834 ] = { 5'd14,	5'd12,	5'd10,	5'd6};
		rom[ 1835 ] = { 5'd2,	5'd7,	5'd18,	5'd9};
		rom[ 1836 ] = { 5'd11,	5'd14,	5'd10,	5'd9};
		rom[ 1837 ] = { 5'd7,	5'd6,	5'd10,	5'd8};
		rom[ 1838 ] = { 5'd6,	5'd6,	5'd14,	5'd6};
		rom[ 1839 ] = { 5'd4,	5'd13,	5'd9,	5'd7};
		rom[ 1840 ] = { 5'd14,	5'd10,	5'd6,	5'd12};
		rom[ 1841 ] = { 5'd4,	5'd10,	5'd6,	5'd12};
		rom[ 1842 ] = { 5'd13,	5'd9,	5'd8,	5'd6};
		rom[ 1843 ] = { 5'd8,	5'd3,	5'd4,	5'd14};
		rom[ 1844 ] = { 5'd17,	5'd0,	5'd3,	5'd18};
		rom[ 1845 ] = { 5'd4,	5'd12,	5'd16,	5'd12};
		rom[ 1846 ] = { 5'd15,	5'd0,	5'd6,	5'd14};
		rom[ 1847 ] = { 5'd3,	5'd0,	5'd6,	5'd14};
		rom[ 1848 ] = { 5'd12,	5'd2,	5'd12,	5'd20};
		rom[ 1849 ] = { 5'd0,	5'd2,	5'd12,	5'd20};
		rom[ 1850 ] = { 5'd16,	5'd0,	5'd6,	5'd17};
		rom[ 1851 ] = { 5'd2,	5'd0,	5'd6,	5'd17};
		rom[ 1852 ] = { 5'd15,	5'd6,	5'd9,	5'd6};
		rom[ 1853 ] = { 5'd0,	5'd6,	5'd9,	5'd6};
		rom[ 1854 ] = { 5'd18,	5'd1,	5'd6,	5'd13};
		rom[ 1855 ] = { 5'd0,	5'd1,	5'd6,	5'd13};
		rom[ 1856 ] = { 5'd16,	5'd0,	5'd4,	5'd9};
		rom[ 1857 ] = { 5'd5,	5'd10,	5'd12,	5'd7};
		rom[ 1858 ] = { 5'd12,	5'd9,	5'd12,	5'd6};
		rom[ 1859 ] = { 5'd0,	5'd9,	5'd12,	5'd6};
		rom[ 1860 ] = { 5'd5,	5'd7,	5'd14,	5'd9};
		rom[ 1861 ] = { 5'd0,	5'd15,	5'd20,	5'd3};
		rom[ 1862 ] = { 5'd8,	5'd10,	5'd8,	5'd10};
		rom[ 1863 ] = { 5'd5,	5'd4,	5'd13,	5'd9};
		rom[ 1864 ] = { 5'd10,	5'd2,	5'd6,	5'd18};
		rom[ 1865 ] = { 5'd6,	5'd0,	5'd6,	5'd9};
		rom[ 1866 ] = { 5'd6,	5'd9,	5'd12,	5'd4};
		rom[ 1867 ] = { 5'd3,	5'd2,	5'd15,	5'd12};
		rom[ 1868 ] = { 5'd12,	5'd0,	5'd12,	5'd5};
		rom[ 1869 ] = { 5'd0,	5'd15,	5'd18,	5'd3};
		rom[ 1870 ] = { 5'd0,	5'd14,	5'd24,	5'd5};
		rom[ 1871 ] = { 5'd5,	5'd1,	5'd3,	5'd18};
		rom[ 1872 ] = { 5'd10,	5'd0,	5'd4,	5'd14};
		rom[ 1873 ] = { 5'd9,	5'd3,	5'd4,	5'd9};
		rom[ 1874 ] = { 5'd8,	5'd2,	5'd12,	5'd6};
		rom[ 1875 ] = { 5'd0,	5'd4,	5'd17,	5'd4};
		rom[ 1876 ] = { 5'd16,	5'd16,	5'd5,	5'd8};
		rom[ 1877 ] = { 5'd3,	5'd16,	5'd5,	5'd8};
		rom[ 1878 ] = { 5'd6,	5'd18,	5'd18,	5'd2};
		rom[ 1879 ] = { 5'd0,	5'd0,	5'd12,	5'd5};
		rom[ 1880 ] = { 5'd14,	5'd3,	5'd6,	5'd12};
		rom[ 1881 ] = { 5'd0,	5'd12,	5'd6,	5'd12};
		rom[ 1882 ] = { 5'd2,	5'd3,	5'd21,	5'd3};
		rom[ 1883 ] = { 5'd4,	5'd3,	5'd6,	5'd12};
		rom[ 1884 ] = { 5'd12,	5'd8,	5'd12,	5'd6};
		rom[ 1885 ] = { 5'd0,	5'd15,	5'd16,	5'd9};
		rom[ 1886 ] = { 5'd6,	5'd13,	5'd18,	5'd5};
		rom[ 1887 ] = { 5'd1,	5'd6,	5'd15,	5'd6};
		rom[ 1888 ] = { 5'd11,	5'd9,	5'd9,	5'd6};
		rom[ 1889 ] = { 5'd3,	5'd0,	5'd15,	5'd11};
		rom[ 1890 ] = { 5'd15,	5'd3,	5'd3,	5'd18};
		rom[ 1891 ] = { 5'd6,	5'd3,	5'd3,	5'd18};
		rom[ 1892 ] = { 5'd9,	5'd5,	5'd10,	5'd8};
		rom[ 1893 ] = { 5'd4,	5'd4,	5'd16,	5'd8};
		rom[ 1894 ] = { 5'd7,	5'd7,	5'd12,	5'd3};
		rom[ 1895 ] = { 5'd5,	5'd0,	5'd9,	5'd13};
		rom[ 1896 ] = { 5'd11,	5'd0,	5'd6,	5'd9};
		rom[ 1897 ] = { 5'd7,	5'd0,	5'd6,	5'd9};
		rom[ 1898 ] = { 5'd8,	5'd1,	5'd10,	5'd9};
		rom[ 1899 ] = { 5'd0,	5'd2,	5'd18,	5'd2};
		rom[ 1900 ] = { 5'd10,	5'd13,	5'd14,	5'd6};
		rom[ 1901 ] = { 5'd0,	5'd13,	5'd14,	5'd6};
		rom[ 1902 ] = { 5'd20,	5'd2,	5'd3,	5'd21};
		rom[ 1903 ] = { 5'd0,	5'd9,	5'd5,	5'd12};
		rom[ 1904 ] = { 5'd12,	5'd6,	5'd12,	5'd6};
		rom[ 1905 ] = { 5'd1,	5'd8,	5'd20,	5'd3};
		rom[ 1906 ] = { 5'd5,	5'd7,	5'd19,	5'd3};
		rom[ 1907 ] = { 5'd1,	5'd12,	5'd9,	5'd6};
		rom[ 1908 ] = { 5'd6,	5'd10,	5'd14,	5'd12};
		rom[ 1909 ] = { 5'd5,	5'd6,	5'd14,	5'd18};
		rom[ 1910 ] = { 5'd11,	5'd12,	5'd9,	5'd7};
		rom[ 1911 ] = { 5'd1,	5'd15,	5'd18,	5'd4};
		rom[ 1912 ] = { 5'd11,	5'd14,	5'd6,	5'd9};
		rom[ 1913 ] = { 5'd0,	5'd8,	5'd18,	5'd4};
		rom[ 1914 ] = { 5'd3,	5'd10,	5'd20,	5'd6};
		rom[ 1915 ] = { 5'd1,	5'd10,	5'd20,	5'd6};
		rom[ 1916 ] = { 5'd0,	5'd9,	5'd24,	5'd2};
		rom[ 1917 ] = { 5'd1,	5'd12,	5'd20,	5'd8};
		rom[ 1918 ] = { 5'd11,	5'd12,	5'd9,	5'd7};
		rom[ 1919 ] = { 5'd4,	5'd12,	5'd9,	5'd7};
		rom[ 1920 ] = { 5'd12,	5'd12,	5'd8,	5'd5};
		rom[ 1921 ] = { 5'd4,	5'd12,	5'd8,	5'd5};
		rom[ 1922 ] = { 5'd13,	5'd10,	5'd4,	5'd10};
		rom[ 1923 ] = { 5'd1,	5'd15,	5'd20,	5'd2};
		rom[ 1924 ] = { 5'd9,	5'd10,	5'd6,	5'd6};
		rom[ 1925 ] = { 5'd0,	5'd1,	5'd21,	5'd3};
		rom[ 1926 ] = { 5'd6,	5'd4,	5'd13,	5'd9};
		rom[ 1927 ] = { 5'd6,	5'd5,	5'd12,	5'd5};
		rom[ 1928 ] = { 5'd10,	5'd10,	5'd10,	5'd6};
		rom[ 1929 ] = { 5'd6,	5'd12,	5'd5,	5'd8};
		rom[ 1930 ] = { 5'd13,	5'd0,	5'd6,	5'd9};
		rom[ 1931 ] = { 5'd2,	5'd10,	5'd18,	5'd6};
		rom[ 1932 ] = { 5'd11,	5'd2,	5'd9,	5'd4};
		rom[ 1933 ] = { 5'd1,	5'd20,	5'd21,	5'd3};
		rom[ 1934 ] = { 5'd1,	5'd10,	5'd22,	5'd2};
		rom[ 1935 ] = { 5'd0,	5'd17,	5'd18,	5'd3};
		rom[ 1936 ] = { 5'd13,	5'd0,	5'd6,	5'd9};
		rom[ 1937 ] = { 5'd5,	5'd0,	5'd6,	5'd9};
		rom[ 1938 ] = { 5'd18,	5'd2,	5'd6,	5'd20};
		rom[ 1939 ] = { 5'd0,	5'd2,	5'd6,	5'd20};
		rom[ 1940 ] = { 5'd11,	5'd7,	5'd6,	5'd14};
		rom[ 1941 ] = { 5'd0,	5'd1,	5'd4,	5'd9};
		rom[ 1942 ] = { 5'd12,	5'd14,	5'd9,	5'd4};
		rom[ 1943 ] = { 5'd1,	5'd13,	5'd9,	5'd4};
		rom[ 1944 ] = { 5'd7,	5'd6,	5'd15,	5'd6};
		rom[ 1945 ] = { 5'd8,	5'd2,	5'd3,	5'd18};
		rom[ 1946 ] = { 5'd6,	5'd6,	5'd12,	5'd6};
		rom[ 1947 ] = { 5'd2,	5'd19,	5'd20,	5'd4};
		rom[ 1948 ] = { 5'd14,	5'd15,	5'd6,	5'd9};
		rom[ 1949 ] = { 5'd3,	5'd5,	5'd18,	5'd14};
		rom[ 1950 ] = { 5'd15,	5'd6,	5'd4,	5'd18};
		rom[ 1951 ] = { 5'd5,	5'd6,	5'd4,	5'd18};
		rom[ 1952 ] = { 5'd11,	5'd0,	5'd6,	5'd9};
		rom[ 1953 ] = { 5'd7,	5'd0,	5'd6,	5'd9};
		rom[ 1954 ] = { 5'd11,	5'd5,	5'd6,	5'd9};
		rom[ 1955 ] = { 5'd9,	5'd5,	5'd6,	5'd6};
		rom[ 1956 ] = { 5'd4,	5'd1,	5'd16,	5'd6};
		rom[ 1957 ] = { 5'd9,	5'd13,	5'd6,	5'd11};
		rom[ 1958 ] = { 5'd17,	5'd1,	5'd6,	5'd12};
		rom[ 1959 ] = { 5'd1,	5'd17,	5'd18,	5'd3};
		rom[ 1960 ] = { 5'd7,	5'd13,	5'd10,	5'd8};
		rom[ 1961 ] = { 5'd6,	5'd18,	5'd10,	5'd6};
		rom[ 1962 ] = { 5'd9,	5'd14,	5'd9,	5'd4};
		rom[ 1963 ] = { 5'd1,	5'd1,	5'd6,	5'd12};
		rom[ 1964 ] = { 5'd19,	5'd4,	5'd5,	5'd12};
		rom[ 1965 ] = { 5'd0,	5'd0,	5'd8,	5'd8};
		rom[ 1966 ] = { 5'd3,	5'd5,	5'd19,	5'd3};
		rom[ 1967 ] = { 5'd1,	5'd5,	5'd12,	5'd6};
		rom[ 1968 ] = { 5'd2,	5'd1,	5'd21,	5'd8};
		rom[ 1969 ] = { 5'd4,	5'd1,	5'd16,	5'd8};
		rom[ 1970 ] = { 5'd6,	5'd0,	5'd18,	5'd3};
		rom[ 1971 ] = { 5'd4,	5'd4,	5'd10,	5'd14};
		rom[ 1972 ] = { 5'd15,	5'd6,	5'd4,	5'd10};
		rom[ 1973 ] = { 5'd3,	5'd18,	5'd18,	5'd3};
		rom[ 1974 ] = { 5'd8,	5'd18,	5'd12,	5'd6};
		rom[ 1975 ] = { 5'd3,	5'd15,	5'd6,	5'd9};
		rom[ 1976 ] = { 5'd15,	5'd7,	5'd6,	5'd8};
		rom[ 1977 ] = { 5'd3,	5'd7,	5'd6,	5'd8};
		rom[ 1978 ] = { 5'd5,	5'd9,	5'd18,	5'd6};
		rom[ 1979 ] = { 5'd1,	5'd13,	5'd12,	5'd6};
		rom[ 1980 ] = { 5'd14,	5'd15,	5'd10,	5'd6};
		rom[ 1981 ] = { 5'd0,	5'd15,	5'd10,	5'd6};
		rom[ 1982 ] = { 5'd15,	5'd13,	5'd6,	5'd9};
		rom[ 1983 ] = { 5'd3,	5'd13,	5'd6,	5'd9};
		rom[ 1984 ] = { 5'd9,	5'd5,	5'd8,	5'd8};
		rom[ 1985 ] = { 5'd1,	5'd18,	5'd12,	5'd6};
		rom[ 1986 ] = { 5'd13,	5'd19,	5'd10,	5'd4};
		rom[ 1987 ] = { 5'd1,	5'd19,	5'd10,	5'd4};
		rom[ 1988 ] = { 5'd6,	5'd19,	5'd18,	5'd3};
		rom[ 1989 ] = { 5'd8,	5'd14,	5'd4,	5'd10};
		rom[ 1990 ] = { 5'd0,	5'd0,	5'd24,	5'd6};
		rom[ 1991 ] = { 5'd0,	5'd1,	5'd6,	5'd9};
		rom[ 1992 ] = { 5'd4,	5'd9,	5'd20,	5'd6};
		rom[ 1993 ] = { 5'd1,	5'd15,	5'd19,	5'd8};
		rom[ 1994 ] = { 5'd14,	5'd0,	5'd10,	5'd6};
		rom[ 1995 ] = { 5'd1,	5'd10,	5'd21,	5'd14};
		rom[ 1996 ] = { 5'd10,	5'd10,	5'd8,	5'd8};
		rom[ 1997 ] = { 5'd6,	5'd8,	5'd10,	5'd4};
		rom[ 1998 ] = { 5'd10,	5'd5,	5'd4,	5'd9};
		rom[ 1999 ] = { 5'd7,	5'd5,	5'd6,	5'd10};
		rom[ 2000 ] = { 5'd14,	5'd4,	5'd4,	5'd13};
		rom[ 2001 ] = { 5'd6,	5'd4,	5'd4,	5'd13};
		rom[ 2002 ] = { 5'd8,	5'd7,	5'd9,	5'd6};
		rom[ 2003 ] = { 5'd3,	5'd6,	5'd16,	5'd6};
		rom[ 2004 ] = { 5'd5,	5'd4,	5'd16,	5'd14};
		rom[ 2005 ] = { 5'd0,	5'd0,	5'd24,	5'd4};
		rom[ 2006 ] = { 5'd9,	5'd1,	5'd9,	5'd6};
		rom[ 2007 ] = { 5'd4,	5'd1,	5'd14,	5'd4};
		rom[ 2008 ] = { 5'd10,	5'd14,	5'd7,	5'd9};
		rom[ 2009 ] = { 5'd8,	5'd3,	5'd8,	5'd10};
		rom[ 2010 ] = { 5'd7,	5'd3,	5'd12,	5'd5};
		rom[ 2011 ] = { 5'd8,	5'd2,	5'd4,	5'd13};
		rom[ 2012 ] = { 5'd11,	5'd2,	5'd3,	5'd19};
		rom[ 2013 ] = { 5'd7,	5'd7,	5'd9,	5'd6};
		rom[ 2014 ] = { 5'd4,	5'd22,	5'd20,	5'd2};
		rom[ 2015 ] = { 5'd0,	5'd16,	5'd24,	5'd4};
		rom[ 2016 ] = { 5'd7,	5'd3,	5'd12,	5'd5};
		rom[ 2017 ] = { 5'd1,	5'd10,	5'd8,	5'd14};
		rom[ 2018 ] = { 5'd11,	5'd16,	5'd6,	5'd6};
		rom[ 2019 ] = { 5'd6,	5'd0,	5'd10,	5'd24};
		rom[ 2020 ] = { 5'd7,	5'd5,	5'd14,	5'd14};
		rom[ 2021 ] = { 5'd7,	5'd8,	5'd10,	5'd8};
		rom[ 2022 ] = { 5'd9,	5'd1,	5'd9,	5'd6};
		rom[ 2023 ] = { 5'd0,	5'd6,	5'd24,	5'd3};
		rom[ 2024 ] = { 5'd7,	5'd3,	5'd12,	5'd5};
		rom[ 2025 ] = { 5'd1,	5'd13,	5'd22,	5'd4};
		rom[ 2026 ] = { 5'd9,	5'd12,	5'd12,	5'd6};
		rom[ 2027 ] = { 5'd0,	5'd5,	5'd9,	5'd6};
		rom[ 2028 ] = { 5'd1,	5'd5,	5'd23,	5'd6};
		rom[ 2029 ] = { 5'd1,	5'd6,	5'd19,	5'd12};
		rom[ 2030 ] = { 5'd9,	5'd1,	5'd6,	5'd21};
		rom[ 2031 ] = { 5'd3,	5'd19,	5'd18,	5'd3};
		rom[ 2032 ] = { 5'd9,	5'd14,	5'd6,	5'd9};
		rom[ 2033 ] = { 5'd9,	5'd6,	5'd4,	5'd12};
		rom[ 2034 ] = { 5'd16,	5'd0,	5'd6,	5'd9};
		rom[ 2035 ] = { 5'd2,	5'd0,	5'd6,	5'd9};
		rom[ 2036 ] = { 5'd13,	5'd1,	5'd4,	5'd22};
		rom[ 2037 ] = { 5'd1,	5'd8,	5'd8,	5'd12};
		rom[ 2038 ] = { 5'd14,	5'd7,	5'd7,	5'd9};
		rom[ 2039 ] = { 5'd3,	5'd12,	5'd18,	5'd4};
		rom[ 2040 ] = { 5'd13,	5'd1,	5'd4,	5'd22};
		rom[ 2041 ] = { 5'd7,	5'd1,	5'd4,	5'd22};
		rom[ 2042 ] = { 5'd4,	5'd7,	5'd20,	5'd4};
		rom[ 2043 ] = { 5'd9,	5'd10,	5'd6,	5'd7};
		rom[ 2044 ] = { 5'd7,	5'd7,	5'd10,	5'd4};
		rom[ 2045 ] = { 5'd0,	5'd3,	5'd4,	5'd15};
		rom[ 2046 ] = { 5'd15,	5'd0,	5'd8,	5'd12};
		rom[ 2047 ] = { 5'd1,	5'd0,	5'd8,	5'd12};
		rom[ 2048 ] = { 5'd14,	5'd5,	5'd6,	5'd16};
		rom[ 2049 ] = { 5'd4,	5'd5,	5'd6,	5'd16};
		rom[ 2050 ] = { 5'd15,	5'd0,	5'd6,	5'd16};
		rom[ 2051 ] = { 5'd3,	5'd0,	5'd6,	5'd16};
		rom[ 2052 ] = { 5'd0,	5'd2,	5'd24,	5'd3};
		rom[ 2053 ] = { 5'd7,	5'd1,	5'd10,	5'd4};
		rom[ 2054 ] = { 5'd1,	5'd0,	5'd23,	5'd8};
		rom[ 2055 ] = { 5'd1,	5'd17,	5'd19,	5'd3};
		rom[ 2056 ] = { 5'd6,	5'd18,	5'd18,	5'd2};
		rom[ 2057 ] = { 5'd1,	5'd17,	5'd9,	5'd6};
		rom[ 2058 ] = { 5'd15,	5'd15,	5'd6,	5'd9};
		rom[ 2059 ] = { 5'd3,	5'd15,	5'd6,	5'd9};
		rom[ 2060 ] = { 5'd4,	5'd14,	5'd20,	5'd6};
		rom[ 2061 ] = { 5'd0,	5'd10,	5'd6,	5'd14};
		rom[ 2062 ] = { 5'd6,	5'd18,	5'd18,	5'd3};
		rom[ 2063 ] = { 5'd4,	5'd12,	5'd9,	5'd7};
		rom[ 2064 ] = { 5'd6,	5'd10,	5'd18,	5'd5};
		rom[ 2065 ] = { 5'd0,	5'd10,	5'd18,	5'd5};
		rom[ 2066 ] = { 5'd3,	5'd2,	5'd18,	5'd9};
		rom[ 2067 ] = { 5'd4,	5'd6,	5'd10,	5'd10};
		rom[ 2068 ] = { 5'd20,	5'd14,	5'd4,	5'd9};
		rom[ 2069 ] = { 5'd0,	5'd14,	5'd4,	5'd9};
		rom[ 2070 ] = { 5'd11,	5'd1,	5'd4,	5'd20};
		rom[ 2071 ] = { 5'd6,	5'd21,	5'd12,	5'd3};
		rom[ 2072 ] = { 5'd11,	5'd1,	5'd4,	5'd20};
		rom[ 2073 ] = { 5'd1,	5'd16,	5'd10,	5'd8};
		rom[ 2074 ] = { 5'd11,	5'd1,	5'd4,	5'd20};
		rom[ 2075 ] = { 5'd1,	5'd0,	5'd3,	5'd19};
		rom[ 2076 ] = { 5'd11,	5'd1,	5'd4,	5'd20};
		rom[ 2077 ] = { 5'd0,	5'd1,	5'd6,	5'd9};
		rom[ 2078 ] = { 5'd3,	5'd7,	5'd19,	5'd4};
		rom[ 2079 ] = { 5'd7,	5'd14,	5'd9,	5'd6};
		rom[ 2080 ] = { 5'd17,	5'd1,	5'd7,	5'd6};
		rom[ 2081 ] = { 5'd5,	5'd0,	5'd14,	5'd8};
		rom[ 2082 ] = { 5'd16,	5'd1,	5'd8,	5'd6};
		rom[ 2083 ] = { 5'd0,	5'd1,	5'd8,	5'd6};
		rom[ 2084 ] = { 5'd6,	5'd0,	5'd18,	5'd4};
		rom[ 2085 ] = { 5'd0,	5'd14,	5'd9,	5'd6};
		rom[ 2086 ] = { 5'd3,	5'd7,	5'd18,	5'd8};
		rom[ 2087 ] = { 5'd2,	5'd11,	5'd6,	5'd9};
		rom[ 2088 ] = { 5'd10,	5'd5,	5'd6,	5'd9};
		rom[ 2089 ] = { 5'd10,	5'd6,	5'd4,	5'd18};
		rom[ 2090 ] = { 5'd11,	5'd1,	5'd4,	5'd20};
		rom[ 2091 ] = { 5'd9,	5'd1,	5'd4,	5'd20};
		rom[ 2092 ] = { 5'd5,	5'd9,	5'd18,	5'd6};
		rom[ 2093 ] = { 5'd6,	5'd4,	5'd6,	5'd9};
		rom[ 2094 ] = { 5'd10,	5'd16,	5'd8,	5'd6};
		rom[ 2095 ] = { 5'd0,	5'd0,	5'd18,	5'd8};
		rom[ 2096 ] = { 5'd6,	5'd5,	5'd14,	5'd12};
		rom[ 2097 ] = { 5'd4,	5'd3,	5'd15,	5'd7};
		rom[ 2098 ] = { 5'd14,	5'd12,	5'd10,	5'd6};
		rom[ 2099 ] = { 5'd0,	5'd11,	5'd4,	5'd10};
		rom[ 2100 ] = { 5'd1,	5'd10,	5'd22,	5'd3};
		rom[ 2101 ] = { 5'd8,	5'd9,	5'd6,	5'd10};
		rom[ 2102 ] = { 5'd13,	5'd2,	5'd6,	5'd12};
		rom[ 2103 ] = { 5'd10,	5'd6,	5'd4,	5'd18};
		rom[ 2104 ] = { 5'd7,	5'd8,	5'd10,	5'd16};
		rom[ 2105 ] = { 5'd8,	5'd1,	5'd8,	5'd12};
		rom[ 2106 ] = { 5'd7,	5'd1,	5'd12,	5'd14};
		rom[ 2107 ] = { 5'd2,	5'd14,	5'd12,	5'd6};
		rom[ 2108 ] = { 5'd11,	5'd16,	5'd6,	5'd6};
		rom[ 2109 ] = { 5'd7,	5'd16,	5'd6,	5'd6};
		rom[ 2110 ] = { 5'd13,	5'd4,	5'd4,	5'd10};
		rom[ 2111 ] = { 5'd0,	5'd19,	5'd19,	5'd3};
		rom[ 2112 ] = { 5'd12,	5'd8,	5'd6,	5'd8};
		rom[ 2113 ] = { 5'd8,	5'd1,	5'd8,	5'd22};
		rom[ 2114 ] = { 5'd12,	5'd8,	5'd6,	5'd8};
		rom[ 2115 ] = { 5'd6,	5'd8,	5'd6,	5'd8};
		rom[ 2116 ] = { 5'd14,	5'd5,	5'd6,	5'd9};
		rom[ 2117 ] = { 5'd0,	5'd6,	5'd24,	5'd4};
		rom[ 2118 ] = { 5'd14,	5'd12,	5'd10,	5'd6};
		rom[ 2119 ] = { 5'd0,	5'd12,	5'd10,	5'd6};
		rom[ 2120 ] = { 5'd4,	5'd6,	5'd19,	5'd3};
		rom[ 2121 ] = { 5'd1,	5'd6,	5'd19,	5'd3};
		rom[ 2122 ] = { 5'd4,	5'd0,	5'd16,	5'd9};
		rom[ 2123 ] = { 5'd0,	5'd1,	5'd24,	5'd5};
		rom[ 2124 ] = { 5'd3,	5'd6,	5'd6,	5'd15};
		rom[ 2125 ] = { 5'd9,	5'd6,	5'd6,	5'd9};
		rom[ 2126 ] = { 5'd0,	5'd17,	5'd18,	5'd3};
		rom[ 2127 ] = { 5'd6,	5'd22,	5'd18,	5'd2};
		rom[ 2128 ] = { 5'd2,	5'd12,	5'd6,	5'd9};
		rom[ 2129 ] = { 5'd18,	5'd12,	5'd6,	5'd9};
		rom[ 2130 ] = { 5'd0,	5'd12,	5'd6,	5'd9};
		rom[ 2131 ] = { 5'd11,	5'd14,	5'd4,	5'd10};
		rom[ 2132 ] = { 5'd9,	5'd6,	5'd6,	5'd16};
		rom[ 2133 ] = { 5'd7,	5'd7,	5'd10,	5'd10};
		rom[ 2134 ] = { 5'd1,	5'd3,	5'd6,	5'd13};
		rom[ 2135 ] = { 5'd18,	5'd1,	5'd6,	5'd13};
		rom[ 2136 ] = { 5'd5,	5'd1,	5'd6,	5'd9};
		rom[ 2137 ] = { 5'd18,	5'd2,	5'd6,	5'd11};
		rom[ 2138 ] = { 5'd0,	5'd2,	5'd6,	5'd11};
		rom[ 2139 ] = { 5'd9,	5'd12,	5'd15,	5'd6};
		rom[ 2140 ] = { 5'd2,	5'd2,	5'd20,	5'd3};
		rom[ 2141 ] = { 5'd10,	5'd6,	5'd4,	5'd9};
		rom[ 2142 ] = { 5'd5,	5'd6,	5'd12,	5'd14};
		rom[ 2143 ] = { 5'd9,	5'd0,	5'd6,	5'd9};
		rom[ 2144 ] = { 5'd7,	5'd0,	5'd9,	5'd6};
		rom[ 2145 ] = { 5'd10,	5'd6,	5'd6,	5'd9};
		rom[ 2146 ] = { 5'd4,	5'd1,	5'd12,	5'd20};
		rom[ 2147 ] = { 5'd6,	5'd7,	5'd18,	5'd3};
		rom[ 2148 ] = { 5'd0,	5'd7,	5'd18,	5'd3};
		rom[ 2149 ] = { 5'd3,	5'd20,	5'd18,	5'd3};
		rom[ 2150 ] = { 5'd9,	5'd6,	5'd6,	5'd9};
		rom[ 2151 ] = { 5'd6,	5'd2,	5'd12,	5'd15};
		rom[ 2152 ] = { 5'd2,	5'd3,	5'd18,	5'd3};
		rom[ 2153 ] = { 5'd19,	5'd4,	5'd4,	5'd18};
		rom[ 2154 ] = { 5'd0,	5'd1,	5'd19,	5'd3};
		rom[ 2155 ] = { 5'd5,	5'd0,	5'd15,	5'd4};
		rom[ 2156 ] = { 5'd5,	5'd2,	5'd14,	5'd5};
		rom[ 2157 ] = { 5'd1,	5'd2,	5'd22,	5'd14};
		rom[ 2158 ] = { 5'd8,	5'd15,	5'd6,	5'd9};
		rom[ 2159 ] = { 5'd6,	5'd17,	5'd18,	5'd3};
		rom[ 2160 ] = { 5'd9,	5'd6,	5'd3,	5'd18};
		rom[ 2161 ] = { 5'd2,	5'd0,	5'd20,	5'd3};
		rom[ 2162 ] = { 5'd5,	5'd4,	5'd5,	5'd12};
		rom[ 2163 ] = { 5'd8,	5'd6,	5'd12,	5'd5};
		rom[ 2164 ] = { 5'd9,	5'd12,	5'd6,	5'd12};
		rom[ 2165 ] = { 5'd14,	5'd14,	5'd8,	5'd10};
		rom[ 2166 ] = { 5'd2,	5'd14,	5'd8,	5'd10};
		rom[ 2167 ] = { 5'd10,	5'd18,	5'd12,	5'd6};
		rom[ 2168 ] = { 5'd1,	5'd3,	5'd6,	5'd9};
		rom[ 2169 ] = { 5'd11,	5'd3,	5'd3,	5'd20};
		rom[ 2170 ] = { 5'd4,	5'd6,	5'd14,	5'd6};
		rom[ 2171 ] = { 5'd6,	5'd5,	5'd12,	5'd13};
		rom[ 2172 ] = { 5'd5,	5'd4,	5'd4,	5'd15};
		rom[ 2173 ] = { 5'd9,	5'd16,	5'd15,	5'd4};
		rom[ 2174 ] = { 5'd7,	5'd8,	5'd6,	5'd14};
		rom[ 2175 ] = { 5'd7,	5'd6,	5'd10,	5'd6};
		rom[ 2176 ] = { 5'd2,	5'd5,	5'd18,	5'd3};
		rom[ 2177 ] = { 5'd5,	5'd1,	5'd15,	5'd8};
		rom[ 2178 ] = { 5'd7,	5'd1,	5'd8,	5'd18};
		rom[ 2179 ] = { 5'd0,	5'd10,	5'd24,	5'd3};
		rom[ 2180 ] = { 5'd0,	5'd2,	5'd6,	5'd13};
		rom[ 2181 ] = { 5'd16,	5'd0,	5'd8,	5'd10};
		rom[ 2182 ] = { 5'd5,	5'd1,	5'd10,	5'd9};
		rom[ 2183 ] = { 5'd5,	5'd6,	5'd18,	5'd3};
		rom[ 2184 ] = { 5'd0,	5'd1,	5'd24,	5'd3};
		rom[ 2185 ] = { 5'd11,	5'd4,	5'd6,	5'd11};
		rom[ 2186 ] = { 5'd0,	5'd0,	5'd8,	5'd10};
		rom[ 2187 ] = { 5'd4,	5'd16,	5'd18,	5'd3};
		rom[ 2188 ] = { 5'd2,	5'd16,	5'd18,	5'd3};
		rom[ 2189 ] = { 5'd3,	5'd0,	5'd18,	5'd10};
		rom[ 2190 ] = { 5'd2,	5'd3,	5'd20,	5'd21};
		rom[ 2191 ] = { 5'd6,	5'd7,	5'd14,	5'd3};
		rom[ 2192 ] = { 5'd0,	5'd9,	5'd12,	5'd6};
		rom[ 2193 ] = { 5'd3,	5'd14,	5'd21,	5'd4};
		rom[ 2194 ] = { 5'd0,	5'd14,	5'd21,	5'd4};
		rom[ 2195 ] = { 5'd5,	5'd21,	5'd18,	5'd3};
		rom[ 2196 ] = { 5'd1,	5'd21,	5'd18,	5'd3};
		rom[ 2197 ] = { 5'd19,	5'd4,	5'd4,	5'd18};
		rom[ 2198 ] = { 5'd3,	5'd7,	5'd18,	5'd3};
		rom[ 2199 ] = { 5'd19,	5'd4,	5'd4,	5'd18};
		rom[ 2200 ] = { 5'd7,	5'd15,	5'd10,	5'd6};
		rom[ 2201 ] = { 5'd9,	5'd13,	5'd11,	5'd9};
		rom[ 2202 ] = { 5'd0,	5'd6,	5'd4,	5'd10};
		rom[ 2203 ] = { 5'd15,	5'd16,	5'd9,	5'd6};
		rom[ 2204 ] = { 5'd1,	5'd5,	5'd4,	5'd18};
		rom[ 2205 ] = { 5'd9,	5'd8,	5'd8,	5'd10};
		rom[ 2206 ] = { 5'd7,	5'd8,	5'd8,	5'd10};
		rom[ 2207 ] = { 5'd9,	5'd8,	5'd12,	5'd5};
		rom[ 2208 ] = { 5'd7,	5'd8,	5'd9,	5'd7};
		rom[ 2209 ] = { 5'd9,	5'd8,	5'd12,	5'd5};
		rom[ 2210 ] = { 5'd7,	5'd6,	5'd9,	5'd7};
		rom[ 2211 ] = { 5'd9,	5'd8,	5'd12,	5'd5};
		rom[ 2212 ] = { 5'd10,	5'd5,	5'd4,	5'd18};
		rom[ 2213 ] = { 5'd5,	5'd5,	5'd14,	5'd12};
		rom[ 2214 ] = { 5'd0,	5'd1,	5'd11,	5'd4};
		rom[ 2215 ] = { 5'd9,	5'd10,	5'd6,	5'd10};
		rom[ 2216 ] = { 5'd2,	5'd17,	5'd11,	5'd6};
		rom[ 2217 ] = { 5'd15,	5'd16,	5'd9,	5'd6};
		rom[ 2218 ] = { 5'd1,	5'd10,	5'd18,	5'd2};
		rom[ 2219 ] = { 5'd6,	5'd4,	5'd12,	5'd13};
		rom[ 2220 ] = { 5'd0,	5'd18,	5'd18,	5'd3};
		rom[ 2221 ] = { 5'd6,	5'd18,	5'd18,	5'd3};
		rom[ 2222 ] = { 5'd0,	5'd16,	5'd9,	5'd6};
		rom[ 2223 ] = { 5'd13,	5'd15,	5'd9,	5'd6};
		rom[ 2224 ] = { 5'd2,	5'd15,	5'd9,	5'd6};
		rom[ 2225 ] = { 5'd13,	5'd1,	5'd6,	5'd16};
		rom[ 2226 ] = { 5'd5,	5'd1,	5'd6,	5'd16};
		rom[ 2227 ] = { 5'd11,	5'd5,	5'd6,	5'd10};
		rom[ 2228 ] = { 5'd7,	5'd5,	5'd6,	5'd10};
		rom[ 2229 ] = { 5'd10,	5'd0,	5'd6,	5'd24};
		rom[ 2230 ] = { 5'd3,	5'd4,	5'd4,	5'd20};
		rom[ 2231 ] = { 5'd14,	5'd0,	5'd6,	5'd9};
		rom[ 2232 ] = { 5'd4,	5'd0,	5'd6,	5'd9};
		rom[ 2233 ] = { 5'd4,	5'd5,	5'd18,	5'd5};
		rom[ 2234 ] = { 5'd5,	5'd6,	5'd6,	5'd9};
		rom[ 2235 ] = { 5'd7,	5'd2,	5'd15,	5'd8};
		rom[ 2236 ] = { 5'd2,	5'd2,	5'd15,	5'd8};
		rom[ 2237 ] = { 5'd10,	5'd0,	5'd4,	5'd9};
		rom[ 2238 ] = { 5'd3,	5'd4,	5'd6,	5'd12};
		rom[ 2239 ] = { 5'd16,	5'd0,	5'd8,	5'd18};
		rom[ 2240 ] = { 5'd0,	5'd0,	5'd8,	5'd18};
		rom[ 2241 ] = { 5'd0,	5'd7,	5'd24,	5'd6};
		rom[ 2242 ] = { 5'd4,	5'd7,	5'd14,	5'd3};
		rom[ 2243 ] = { 5'd10,	5'd8,	5'd8,	5'd15};
		rom[ 2244 ] = { 5'd7,	5'd0,	5'd10,	5'd14};
		rom[ 2245 ] = { 5'd13,	5'd10,	5'd8,	5'd10};
		rom[ 2246 ] = { 5'd3,	5'd0,	5'd4,	5'd9};
		rom[ 2247 ] = { 5'd16,	5'd1,	5'd6,	5'd8};
		rom[ 2248 ] = { 5'd2,	5'd1,	5'd6,	5'd8};
		rom[ 2249 ] = { 5'd3,	5'd6,	5'd18,	5'd12};
		rom[ 2250 ] = { 5'd4,	5'd12,	5'd16,	5'd4};
		rom[ 2251 ] = { 5'd4,	5'd9,	5'd16,	5'd15};
		rom[ 2252 ] = { 5'd3,	5'd10,	5'd8,	5'd10};
		rom[ 2253 ] = { 5'd8,	5'd18,	5'd16,	5'd6};
		rom[ 2254 ] = { 5'd2,	5'd16,	5'd12,	5'd5};
		rom[ 2255 ] = { 5'd14,	5'd14,	5'd9,	5'd4};
		rom[ 2256 ] = { 5'd7,	5'd14,	5'd9,	5'd6};
		rom[ 2257 ] = { 5'd4,	5'd10,	5'd16,	5'd12};
		rom[ 2258 ] = { 5'd0,	5'd13,	5'd19,	5'd6};
		rom[ 2259 ] = { 5'd10,	5'd13,	5'd9,	5'd6};
		rom[ 2260 ] = { 5'd5,	5'd0,	5'd3,	5'd23};
		rom[ 2261 ] = { 5'd0,	5'd8,	5'd24,	5'd6};
		rom[ 2262 ] = { 5'd0,	5'd5,	5'd5,	5'd12};
		rom[ 2263 ] = { 5'd3,	5'd0,	5'd19,	5'd18};
		rom[ 2264 ] = { 5'd9,	5'd11,	5'd6,	5'd12};
		rom[ 2265 ] = { 5'd0,	5'd5,	5'd24,	5'd8};
		rom[ 2266 ] = { 5'd6,	5'd18,	5'd9,	5'd4};
		rom[ 2267 ] = { 5'd8,	5'd8,	5'd10,	5'd6};
		rom[ 2268 ] = { 5'd2,	5'd7,	5'd20,	5'd3};
		rom[ 2269 ] = { 5'd12,	5'd0,	5'd7,	5'd20};
		rom[ 2270 ] = { 5'd5,	5'd0,	5'd7,	5'd20};
		rom[ 2271 ] = { 5'd14,	5'd2,	5'd2,	5'd18};
		rom[ 2272 ] = { 5'd5,	5'd8,	5'd10,	5'd12};
		rom[ 2273 ] = { 5'd6,	5'd9,	5'd12,	5'd8};
		rom[ 2274 ] = { 5'd7,	5'd7,	5'd3,	5'd14};
		rom[ 2275 ] = { 5'd11,	5'd2,	5'd12,	5'd16};
		rom[ 2276 ] = { 5'd7,	5'd0,	5'd6,	5'd9};
		rom[ 2277 ] = { 5'd13,	5'd14,	5'd9,	5'd4};
		rom[ 2278 ] = { 5'd0,	5'd12,	5'd22,	5'd4};
		rom[ 2279 ] = { 5'd1,	5'd12,	5'd22,	5'd6};
		rom[ 2280 ] = { 5'd6,	5'd6,	5'd9,	5'd6};
		rom[ 2281 ] = { 5'd10,	5'd0,	5'd4,	5'd9};
		rom[ 2282 ] = { 5'd3,	5'd8,	5'd18,	5'd7};
		rom[ 2283 ] = { 5'd0,	5'd6,	5'd24,	5'd6};
		rom[ 2284 ] = { 5'd0,	5'd11,	5'd24,	5'd10};
		rom[ 2285 ] = { 5'd3,	5'd3,	5'd18,	5'd21};
		rom[ 2286 ] = { 5'd7,	5'd12,	5'd4,	5'd10};
		rom[ 2287 ] = { 5'd10,	5'd16,	5'd10,	5'd8};
		rom[ 2288 ] = { 5'd8,	5'd6,	5'd6,	5'd9};
		rom[ 2289 ] = { 5'd12,	5'd10,	5'd6,	5'd12};
		rom[ 2290 ] = { 5'd6,	5'd10,	5'd6,	5'd12};
		rom[ 2291 ] = { 5'd16,	5'd12,	5'd6,	5'd12};
		rom[ 2292 ] = { 5'd2,	5'd12,	5'd6,	5'd12};
		rom[ 2293 ] = { 5'd10,	5'd15,	5'd6,	5'd9};
		rom[ 2294 ] = { 5'd8,	5'd15,	5'd6,	5'd9};
		rom[ 2295 ] = { 5'd14,	5'd20,	5'd10,	5'd4};
		rom[ 2296 ] = { 5'd0,	5'd20,	5'd10,	5'd4};
		rom[ 2297 ] = { 5'd11,	5'd17,	5'd9,	5'd6};
		rom[ 2298 ] = { 5'd3,	5'd2,	5'd14,	5'd4};
		rom[ 2299 ] = { 5'd10,	5'd1,	5'd10,	5'd4};
		rom[ 2300 ] = { 5'd0,	5'd15,	5'd10,	5'd4};
		rom[ 2301 ] = { 5'd19,	5'd2,	5'd3,	5'd19};
		rom[ 2302 ] = { 5'd4,	5'd12,	5'd9,	5'd8};
		rom[ 2303 ] = { 5'd4,	5'd7,	5'd5,	5'd12};
		rom[ 2304 ] = { 5'd0,	5'd1,	5'd24,	5'd3};
		rom[ 2305 ] = { 5'd6,	5'd8,	5'd12,	5'd4};
		rom[ 2306 ] = { 5'd19,	5'd3,	5'd4,	5'd10};
		rom[ 2307 ] = { 5'd0,	5'd6,	5'd9,	5'd6};
		rom[ 2308 ] = { 5'd18,	5'd0,	5'd6,	5'd22};
		rom[ 2309 ] = { 5'd0,	5'd0,	5'd6,	5'd22};
		rom[ 2310 ] = { 5'd5,	5'd15,	5'd19,	5'd3};
		rom[ 2311 ] = { 5'd10,	5'd7,	5'd4,	5'd15};
		rom[ 2312 ] = { 5'd9,	5'd6,	5'd6,	5'd9};
		rom[ 2313 ] = { 5'd0,	5'd21,	5'd18,	5'd3};
		rom[ 2314 ] = { 5'd7,	5'd3,	5'd10,	5'd15};
		rom[ 2315 ] = { 5'd1,	5'd7,	5'd18,	5'd3};
		rom[ 2316 ] = { 5'd8,	5'd2,	5'd9,	5'd6};
		rom[ 2317 ] = { 5'd0,	5'd10,	5'd24,	5'd14};
		rom[ 2318 ] = { 5'd13,	5'd9,	5'd8,	5'd10};
		rom[ 2319 ] = { 5'd10,	5'd5,	5'd4,	5'd9};
		rom[ 2320 ] = { 5'd13,	5'd9,	5'd8,	5'd10};
		rom[ 2321 ] = { 5'd7,	5'd11,	5'd10,	5'd10};
		rom[ 2322 ] = { 5'd4,	5'd13,	5'd18,	5'd4};
		rom[ 2323 ] = { 5'd0,	5'd0,	5'd19,	5'd2};
		rom[ 2324 ] = { 5'd0,	5'd18,	5'd24,	5'd6};
		rom[ 2325 ] = { 5'd6,	5'd4,	5'd8,	5'd16};
		rom[ 2326 ] = { 5'd7,	5'd8,	5'd10,	5'd4};
		rom[ 2327 ] = { 5'd0,	5'd3,	5'd6,	5'd9};
		rom[ 2328 ] = { 5'd13,	5'd15,	5'd7,	5'd9};
		rom[ 2329 ] = { 5'd3,	5'd18,	5'd12,	5'd6};
		rom[ 2330 ] = { 5'd12,	5'd14,	5'd6,	5'd9};
		rom[ 2331 ] = { 5'd2,	5'd15,	5'd15,	5'd8};
		rom[ 2332 ] = { 5'd9,	5'd6,	5'd6,	5'd16};
		rom[ 2333 ] = { 5'd6,	5'd6,	5'd7,	5'd12};
		rom[ 2334 ] = { 5'd14,	5'd6,	5'd6,	5'd9};
		rom[ 2335 ] = { 5'd5,	5'd14,	5'd6,	5'd9};
		rom[ 2336 ] = { 5'd10,	5'd8,	5'd6,	5'd9};
		rom[ 2337 ] = { 5'd6,	5'd6,	5'd4,	5'd18};
		rom[ 2338 ] = { 5'd14,	5'd9,	5'd6,	5'd12};
		rom[ 2339 ] = { 5'd4,	5'd9,	5'd6,	5'd12};
		rom[ 2340 ] = { 5'd14,	5'd15,	5'd9,	5'd6};
		rom[ 2341 ] = { 5'd0,	5'd20,	5'd18,	5'd4};
		rom[ 2342 ] = { 5'd13,	5'd18,	5'd9,	5'd6};
		rom[ 2343 ] = { 5'd2,	5'd18,	5'd9,	5'd6};
		rom[ 2344 ] = { 5'd6,	5'd16,	5'd18,	5'd3};
		rom[ 2345 ] = { 5'd0,	5'd16,	5'd18,	5'd3};
		rom[ 2346 ] = { 5'd19,	5'd2,	5'd4,	5'd22};
		rom[ 2347 ] = { 5'd1,	5'd2,	5'd4,	5'd22};
		rom[ 2348 ] = { 5'd15,	5'd0,	5'd2,	5'd24};
		rom[ 2349 ] = { 5'd3,	5'd20,	5'd16,	5'd4};
		rom[ 2350 ] = { 5'd11,	5'd6,	5'd4,	5'd18};
		rom[ 2351 ] = { 5'd7,	5'd9,	5'd10,	5'd14};
		rom[ 2352 ] = { 5'd14,	5'd6,	5'd6,	5'd9};
		rom[ 2353 ] = { 5'd3,	5'd6,	5'd7,	5'd9};
		rom[ 2354 ] = { 5'd20,	5'd4,	5'd4,	5'd20};
		rom[ 2355 ] = { 5'd7,	5'd6,	5'd6,	5'd9};
		rom[ 2356 ] = { 5'd7,	5'd0,	5'd10,	5'd14};
		rom[ 2357 ] = { 5'd2,	5'd1,	5'd18,	5'd6};
		rom[ 2358 ] = { 5'd15,	5'd0,	5'd2,	5'd24};
		rom[ 2359 ] = { 5'd7,	5'd0,	5'd2,	5'd24};
		rom[ 2360 ] = { 5'd13,	5'd12,	5'd6,	5'd7};
		rom[ 2361 ] = { 5'd5,	5'd12,	5'd6,	5'd7};
		rom[ 2362 ] = { 5'd3,	5'd5,	5'd18,	5'd19};
		rom[ 2363 ] = { 5'd5,	5'd6,	5'd9,	5'd6};
		rom[ 2364 ] = { 5'd9,	5'd5,	5'd9,	5'd6};
		rom[ 2365 ] = { 5'd3,	5'd16,	5'd10,	5'd8};
		rom[ 2366 ] = { 5'd19,	5'd8,	5'd5,	5'd15};
		rom[ 2367 ] = { 5'd0,	5'd8,	5'd5,	5'd15};
		rom[ 2368 ] = { 5'd20,	5'd4,	5'd4,	5'd20};
		rom[ 2369 ] = { 5'd0,	5'd4,	5'd4,	5'd20};
		rom[ 2370 ] = { 5'd7,	5'd7,	5'd10,	5'd4};
		rom[ 2371 ] = { 5'd4,	5'd19,	5'd14,	5'd4};
		rom[ 2372 ] = { 5'd10,	5'd11,	5'd12,	5'd3};
		rom[ 2373 ] = { 5'd0,	5'd1,	5'd24,	5'd3};
		rom[ 2374 ] = { 5'd7,	5'd2,	5'd14,	5'd20};
		rom[ 2375 ] = { 5'd0,	5'd13,	5'd6,	5'd9};
		rom[ 2376 ] = { 5'd13,	5'd0,	5'd4,	5'd19};
		rom[ 2377 ] = { 5'd1,	5'd11,	5'd14,	5'd3};
		rom[ 2378 ] = { 5'd7,	5'd1,	5'd16,	5'd20};
		rom[ 2379 ] = { 5'd0,	5'd10,	5'd21,	5'd9};
		rom[ 2380 ] = { 5'd6,	5'd19,	5'd15,	5'd5};
		rom[ 2381 ] = { 5'd8,	5'd10,	5'd6,	5'd6};
		rom[ 2382 ] = { 5'd7,	5'd1,	5'd16,	5'd20};
		rom[ 2383 ] = { 5'd1,	5'd1,	5'd16,	5'd20};
		rom[ 2384 ] = { 5'd16,	5'd4,	5'd3,	5'd12};
		rom[ 2385 ] = { 5'd5,	5'd4,	5'd3,	5'd12};
		rom[ 2386 ] = { 5'd7,	5'd6,	5'd10,	5'd8};
		rom[ 2387 ] = { 5'd4,	5'd9,	5'd6,	5'd6};
		rom[ 2388 ] = { 5'd6,	5'd5,	5'd12,	5'd4};
		rom[ 2389 ] = { 5'd9,	5'd2,	5'd5,	5'd15};
		rom[ 2390 ] = { 5'd15,	5'd0,	5'd9,	5'd6};
		rom[ 2391 ] = { 5'd6,	5'd0,	5'd11,	5'd10};
		rom[ 2392 ] = { 5'd12,	5'd7,	5'd4,	5'd12};
		rom[ 2393 ] = { 5'd7,	5'd2,	5'd9,	5'd4};
		rom[ 2394 ] = { 5'd6,	5'd0,	5'd13,	5'd6};
		rom[ 2395 ] = { 5'd10,	5'd6,	5'd4,	5'd18};
		rom[ 2396 ] = { 5'd10,	5'd8,	5'd6,	5'd9};
		rom[ 2397 ] = { 5'd3,	5'd18,	5'd10,	5'd6};
		rom[ 2398 ] = { 5'd4,	5'd14,	5'd20,	5'd3};
		rom[ 2399 ] = { 5'd2,	5'd15,	5'd9,	5'd6};
		rom[ 2400 ] = { 5'd13,	5'd0,	5'd4,	5'd19};
		rom[ 2401 ] = { 5'd7,	5'd0,	5'd4,	5'd19};
		rom[ 2402 ] = { 5'd1,	5'd4,	5'd22,	5'd2};
		rom[ 2403 ] = { 5'd0,	5'd0,	5'd9,	5'd6};
		rom[ 2404 ] = { 5'd0,	5'd0,	5'd24,	5'd18};
		rom[ 2405 ] = { 5'd3,	5'd2,	5'd16,	5'd8};
		rom[ 2406 ] = { 5'd3,	5'd6,	5'd18,	5'd6};
		rom[ 2407 ] = { 5'd3,	5'd1,	5'd6,	5'd10};
		rom[ 2408 ] = { 5'd13,	5'd0,	5'd9,	5'd6};
		rom[ 2409 ] = { 5'd2,	5'd0,	5'd9,	5'd6};
		rom[ 2410 ] = { 5'd10,	5'd2,	5'd4,	5'd15};
		rom[ 2411 ] = { 5'd6,	5'd0,	5'd7,	5'd10};
		rom[ 2412 ] = { 5'd2,	5'd2,	5'd20,	5'd4};
		rom[ 2413 ] = { 5'd2,	5'd11,	5'd19,	5'd3};
		rom[ 2414 ] = { 5'd10,	5'd8,	5'd6,	5'd9};
		rom[ 2415 ] = { 5'd8,	5'd8,	5'd6,	5'd9};
		rom[ 2416 ] = { 5'd13,	5'd8,	5'd4,	5'd9};
		rom[ 2417 ] = { 5'd3,	5'd11,	5'd9,	5'd9};
		rom[ 2418 ] = { 5'd3,	5'd9,	5'd18,	5'd5};
		rom[ 2419 ] = { 5'd2,	5'd4,	5'd2,	5'd20};
		rom[ 2420 ] = { 5'd14,	5'd17,	5'd8,	5'd6};
		rom[ 2421 ] = { 5'd3,	5'd21,	5'd18,	5'd2};
		rom[ 2422 ] = { 5'd5,	5'd4,	5'd15,	5'd6};
		rom[ 2423 ] = { 5'd2,	5'd15,	5'd12,	5'd6};
		rom[ 2424 ] = { 5'd17,	5'd8,	5'd6,	5'd9};
		rom[ 2425 ] = { 5'd2,	5'd12,	5'd20,	5'd4};
		rom[ 2426 ] = { 5'd0,	5'd17,	5'd24,	5'd6};
		rom[ 2427 ] = { 5'd7,	5'd16,	5'd9,	5'd4};
		rom[ 2428 ] = { 5'd15,	5'd1,	5'd4,	5'd22};
		rom[ 2429 ] = { 5'd5,	5'd1,	5'd4,	5'd22};
		rom[ 2430 ] = { 5'd11,	5'd13,	5'd8,	5'd9};
		rom[ 2431 ] = { 5'd6,	5'd1,	5'd6,	5'd9};
		rom[ 2432 ] = { 5'd11,	5'd4,	5'd3,	5'd18};
		rom[ 2433 ] = { 5'd5,	5'd8,	5'd12,	5'd6};
		rom[ 2434 ] = { 5'd15,	5'd7,	5'd5,	5'd8};
		rom[ 2435 ] = { 5'd4,	5'd7,	5'd5,	5'd8};
		rom[ 2436 ] = { 5'd12,	5'd6,	5'd6,	5'd12};
		rom[ 2437 ] = { 5'd6,	5'd6,	5'd6,	5'd12};
		rom[ 2438 ] = { 5'd5,	5'd9,	5'd14,	5'd8};
		rom[ 2439 ] = { 5'd9,	5'd1,	5'd3,	5'd14};
		rom[ 2440 ] = { 5'd12,	5'd6,	5'd6,	5'd12};
		rom[ 2441 ] = { 5'd4,	5'd5,	5'd4,	5'd18};
		rom[ 2442 ] = { 5'd4,	5'd6,	5'd16,	5'd18};
		rom[ 2443 ] = { 5'd5,	5'd4,	5'd7,	5'd20};
		rom[ 2444 ] = { 5'd14,	5'd8,	5'd8,	5'd12};
		rom[ 2445 ] = { 5'd9,	5'd10,	5'd6,	5'd14};
		rom[ 2446 ] = { 5'd9,	5'd5,	5'd9,	5'd6};
		rom[ 2447 ] = { 5'd9,	5'd4,	5'd3,	5'd18};
		rom[ 2448 ] = { 5'd1,	5'd4,	5'd22,	5'd14};
		rom[ 2449 ] = { 5'd2,	5'd7,	5'd18,	5'd2};
		rom[ 2450 ] = { 5'd12,	5'd6,	5'd6,	5'd12};
		rom[ 2451 ] = { 5'd6,	5'd5,	5'd9,	5'd7};
		rom[ 2452 ] = { 5'd12,	5'd7,	5'd4,	5'd12};
		rom[ 2453 ] = { 5'd8,	5'd7,	5'd4,	5'd12};
		rom[ 2454 ] = { 5'd7,	5'd2,	5'd10,	5'd22};
		rom[ 2455 ] = { 5'd0,	5'd1,	5'd3,	5'd20};
		rom[ 2456 ] = { 5'd4,	5'd13,	5'd18,	5'd4};
		rom[ 2457 ] = { 5'd2,	5'd13,	5'd18,	5'd4};
		rom[ 2458 ] = { 5'd15,	5'd15,	5'd9,	5'd6};
		rom[ 2459 ] = { 5'd0,	5'd15,	5'd9,	5'd6};
		rom[ 2460 ] = { 5'd6,	5'd0,	5'd18,	5'd24};
		rom[ 2461 ] = { 5'd6,	5'd6,	5'd6,	5'd12};
		rom[ 2462 ] = { 5'd8,	5'd7,	5'd10,	5'd4};
		rom[ 2463 ] = { 5'd1,	5'd9,	5'd18,	5'd6};
		rom[ 2464 ] = { 5'd6,	5'd6,	5'd18,	5'd3};
		rom[ 2465 ] = { 5'd7,	5'd7,	5'd9,	5'd8};
		rom[ 2466 ] = { 5'd10,	5'd12,	5'd6,	5'd12};
		rom[ 2467 ] = { 5'd3,	5'd14,	5'd18,	5'd3};
		rom[ 2468 ] = { 5'd15,	5'd17,	5'd9,	5'd7};
		rom[ 2469 ] = { 5'd1,	5'd12,	5'd10,	5'd6};
		rom[ 2470 ] = { 5'd15,	5'd17,	5'd9,	5'd7};
		rom[ 2471 ] = { 5'd10,	5'd3,	5'd3,	5'd19};
		rom[ 2472 ] = { 5'd15,	5'd17,	5'd9,	5'd7};
		rom[ 2473 ] = { 5'd6,	5'd1,	5'd11,	5'd9};
		rom[ 2474 ] = { 5'd15,	5'd17,	5'd9,	5'd7};
		rom[ 2475 ] = { 5'd6,	5'd5,	5'd11,	5'd6};
		rom[ 2476 ] = { 5'd16,	5'd7,	5'd8,	5'd5};
		rom[ 2477 ] = { 5'd2,	5'd4,	5'd20,	5'd19};
		rom[ 2478 ] = { 5'd2,	5'd1,	5'd21,	5'd6};
		rom[ 2479 ] = { 5'd6,	5'd5,	5'd12,	5'd14};
		rom[ 2480 ] = { 5'd9,	5'd0,	5'd6,	5'd9};
		rom[ 2481 ] = { 5'd2,	5'd11,	5'd8,	5'd5};
		rom[ 2482 ] = { 5'd16,	5'd7,	5'd8,	5'd5};
		rom[ 2483 ] = { 5'd0,	5'd7,	5'd8,	5'd5};
		rom[ 2484 ] = { 5'd15,	5'd17,	5'd9,	5'd7};
		rom[ 2485 ] = { 5'd8,	5'd6,	5'd8,	5'd10};
		rom[ 2486 ] = { 5'd15,	5'd15,	5'd9,	5'd9};
		rom[ 2487 ] = { 5'd0,	5'd15,	5'd9,	5'd9};
		rom[ 2488 ] = { 5'd12,	5'd10,	5'd9,	5'd7};
		rom[ 2489 ] = { 5'd3,	5'd10,	5'd9,	5'd7};
		rom[ 2490 ] = { 5'd13,	5'd15,	5'd10,	5'd8};
		rom[ 2491 ] = { 5'd0,	5'd1,	5'd6,	5'd12};
		rom[ 2492 ] = { 5'd10,	5'd0,	5'd6,	5'd12};
		rom[ 2493 ] = { 5'd7,	5'd0,	5'd10,	5'd12};
		rom[ 2494 ] = { 5'd4,	5'd1,	5'd16,	5'd8};
		rom[ 2495 ] = { 5'd0,	5'd21,	5'd19,	5'd3};
		rom[ 2496 ] = { 5'd6,	5'd9,	5'd18,	5'd4};
		rom[ 2497 ] = { 5'd3,	5'd4,	5'd9,	5'd6};
		rom[ 2498 ] = { 5'd9,	5'd1,	5'd6,	5'd15};
		rom[ 2499 ] = { 5'd5,	5'd9,	5'd6,	5'd6};
		rom[ 2500 ] = { 5'd5,	5'd1,	5'd14,	5'd9};
		rom[ 2501 ] = { 5'd3,	5'd0,	5'd8,	5'd20};
		rom[ 2502 ] = { 5'd5,	5'd0,	5'd7,	5'd9};
		rom[ 2503 ] = { 5'd6,	5'd6,	5'd12,	5'd5};
		rom[ 2504 ] = { 5'd0,	5'd1,	5'd8,	5'd14};
		rom[ 2505 ] = { 5'd2,	5'd12,	5'd22,	5'd4};
		rom[ 2506 ] = { 5'd8,	5'd17,	5'd6,	5'd6};
		rom[ 2507 ] = { 5'd18,	5'd1,	5'd6,	5'd7};
		rom[ 2508 ] = { 5'd0,	5'd0,	5'd6,	5'd6};
		rom[ 2509 ] = { 5'd4,	5'd6,	5'd17,	5'd18};
		rom[ 2510 ] = { 5'd6,	5'd0,	5'd12,	5'd6};
		rom[ 2511 ] = { 5'd4,	5'd7,	5'd18,	5'd4};
		rom[ 2512 ] = { 5'd4,	5'd12,	5'd10,	5'd6};
		rom[ 2513 ] = { 5'd7,	5'd9,	5'd10,	5'd12};
		rom[ 2514 ] = { 5'd0,	5'd1,	5'd24,	5'd3};
		rom[ 2515 ] = { 5'd13,	5'd11,	5'd6,	5'd6};
		rom[ 2516 ] = { 5'd5,	5'd11,	5'd6,	5'd6};
		rom[ 2517 ] = { 5'd3,	5'd10,	5'd19,	5'd3};
		rom[ 2518 ] = { 5'd0,	5'd2,	5'd6,	5'd9};
		rom[ 2519 ] = { 5'd14,	5'd16,	5'd10,	5'd6};
		rom[ 2520 ] = { 5'd0,	5'd16,	5'd10,	5'd6};
		rom[ 2521 ] = { 5'd14,	5'd13,	5'd9,	5'd6};
		rom[ 2522 ] = { 5'd0,	5'd16,	5'd18,	5'd3};
		rom[ 2523 ] = { 5'd6,	5'd16,	5'd18,	5'd3};
		rom[ 2524 ] = { 5'd0,	5'd18,	5'd9,	5'd6};
		rom[ 2525 ] = { 5'd14,	5'd13,	5'd9,	5'd6};
		rom[ 2526 ] = { 5'd6,	5'd2,	5'd6,	5'd9};
		rom[ 2527 ] = { 5'd15,	5'd8,	5'd4,	5'd12};
		rom[ 2528 ] = { 5'd8,	5'd13,	5'd8,	5'd8};
		rom[ 2529 ] = { 5'd4,	5'd20,	5'd18,	5'd3};
		rom[ 2530 ] = { 5'd5,	5'd8,	5'd4,	5'd12};
		rom[ 2531 ] = { 5'd7,	5'd7,	5'd12,	5'd3};
		rom[ 2532 ] = { 5'd10,	5'd6,	5'd4,	5'd9};
		rom[ 2533 ] = { 5'd5,	5'd20,	5'd18,	5'd3};
		rom[ 2534 ] = { 5'd1,	5'd20,	5'd18,	5'd3};
		rom[ 2535 ] = { 5'd18,	5'd1,	5'd6,	5'd20};
		rom[ 2536 ] = { 5'd0,	5'd1,	5'd6,	5'd20};
		rom[ 2537 ] = { 5'd13,	5'd3,	5'd4,	5'd18};
		rom[ 2538 ] = { 5'd0,	5'd2,	5'd6,	5'd12};
		rom[ 2539 ] = { 5'd12,	5'd9,	5'd12,	5'd6};
		rom[ 2540 ] = { 5'd7,	5'd3,	5'd4,	5'd18};
		rom[ 2541 ] = { 5'd14,	5'd0,	5'd6,	5'd9};
		rom[ 2542 ] = { 5'd0,	5'd9,	5'd12,	5'd6};
		rom[ 2543 ] = { 5'd14,	5'd4,	5'd8,	5'd20};
		rom[ 2544 ] = { 5'd2,	5'd4,	5'd8,	5'd20};
		rom[ 2545 ] = { 5'd14,	5'd13,	5'd9,	5'd6};
		rom[ 2546 ] = { 5'd1,	5'd13,	5'd9,	5'd6};
		rom[ 2547 ] = { 5'd3,	5'd15,	5'd18,	5'd3};
		rom[ 2548 ] = { 5'd5,	5'd13,	5'd9,	5'd6};
		rom[ 2549 ] = { 5'd5,	5'd0,	5'd18,	5'd3};
		rom[ 2550 ] = { 5'd8,	5'd2,	5'd6,	5'd7};
		rom[ 2551 ] = { 5'd9,	5'd1,	5'd9,	5'd6};
		rom[ 2552 ] = { 5'd6,	5'd1,	5'd9,	5'd6};
		rom[ 2553 ] = { 5'd5,	5'd6,	5'd14,	5'd6};
		rom[ 2554 ] = { 5'd8,	5'd2,	5'd6,	5'd13};
		rom[ 2555 ] = { 5'd6,	5'd11,	5'd12,	5'd6};
		rom[ 2556 ] = { 5'd3,	5'd1,	5'd18,	5'd15};
		rom[ 2557 ] = { 5'd13,	5'd0,	5'd6,	5'd7};
		rom[ 2558 ] = { 5'd3,	5'd3,	5'd16,	5'd6};
		rom[ 2559 ] = { 5'd12,	5'd1,	5'd3,	5'd12};
		rom[ 2560 ] = { 5'd7,	5'd7,	5'd6,	5'd9};
		rom[ 2561 ] = { 5'd13,	5'd0,	5'd4,	5'd24};
		rom[ 2562 ] = { 5'd7,	5'd0,	5'd4,	5'd24};
		rom[ 2563 ] = { 5'd11,	5'd9,	5'd5,	5'd12};
		rom[ 2564 ] = { 5'd7,	5'd15,	5'd9,	5'd6};
		rom[ 2565 ] = { 5'd5,	5'd7,	5'd18,	5'd6};
		rom[ 2566 ] = { 5'd8,	5'd9,	5'd5,	5'd12};
		rom[ 2567 ] = { 5'd4,	5'd17,	5'd17,	5'd6};
		rom[ 2568 ] = { 5'd0,	5'd3,	5'd18,	5'd14};
		rom[ 2569 ] = { 5'd0,	5'd1,	5'd24,	5'd2};
		rom[ 2570 ] = { 5'd0,	5'd15,	5'd18,	5'd3};
		rom[ 2571 ] = { 5'd9,	5'd0,	5'd6,	5'd9};
		rom[ 2572 ] = { 5'd3,	5'd3,	5'd14,	5'd12};
		rom[ 2573 ] = { 5'd12,	5'd1,	5'd3,	5'd12};
		rom[ 2574 ] = { 5'd8,	5'd0,	5'd6,	5'd9};
		rom[ 2575 ] = { 5'd10,	5'd6,	5'd6,	5'd10};
		rom[ 2576 ] = { 5'd5,	5'd0,	5'd6,	5'd9};
		rom[ 2577 ] = { 5'd2,	5'd0,	5'd21,	5'd7};
		rom[ 2578 ] = { 5'd6,	5'd11,	5'd12,	5'd5};
		rom[ 2579 ] = { 5'd8,	5'd7,	5'd9,	5'd8};
		rom[ 2580 ] = { 5'd9,	5'd6,	5'd6,	5'd18};
		rom[ 2581 ] = { 5'd15,	5'd14,	5'd8,	5'd10};
		rom[ 2582 ] = { 5'd1,	5'd14,	5'd8,	5'd10};
		rom[ 2583 ] = { 5'd11,	5'd0,	5'd8,	5'd10};
		rom[ 2584 ] = { 5'd5,	5'd0,	5'd8,	5'd10};
		rom[ 2585 ] = { 5'd6,	5'd1,	5'd12,	5'd5};
		rom[ 2586 ] = { 5'd1,	5'd12,	5'd18,	5'd2};
		rom[ 2587 ] = { 5'd2,	5'd8,	5'd20,	5'd6};
		rom[ 2588 ] = { 5'd7,	5'd6,	5'd9,	5'd7};
		rom[ 2589 ] = { 5'd10,	5'd5,	5'd8,	5'd16};
		rom[ 2590 ] = { 5'd3,	5'd9,	5'd16,	5'd8};
		rom[ 2591 ] = { 5'd7,	5'd8,	5'd10,	5'd4};
		rom[ 2592 ] = { 5'd7,	5'd12,	5'd10,	5'd8};
		rom[ 2593 ] = { 5'd9,	5'd19,	5'd15,	5'd4};
		rom[ 2594 ] = { 5'd1,	5'd0,	5'd18,	5'd9};
		rom[ 2595 ] = { 5'd13,	5'd4,	5'd10,	5'd8};
		rom[ 2596 ] = { 5'd3,	5'd16,	5'd18,	5'd4};
		rom[ 2597 ] = { 5'd8,	5'd7,	5'd10,	5'd12};
		rom[ 2598 ] = { 5'd6,	5'd7,	5'd10,	5'd12};
		rom[ 2599 ] = { 5'd4,	5'd6,	5'd18,	5'd7};
		rom[ 2600 ] = { 5'd0,	5'd17,	5'd18,	5'd3};
		rom[ 2601 ] = { 5'd3,	5'd17,	5'd18,	5'd3};
		rom[ 2602 ] = { 5'd2,	5'd4,	5'd6,	5'd10};
		rom[ 2603 ] = { 5'd16,	5'd0,	5'd8,	5'd24};
		rom[ 2604 ] = { 5'd4,	5'd0,	5'd8,	5'd15};
		rom[ 2605 ] = { 5'd16,	5'd0,	5'd8,	5'd24};
		rom[ 2606 ] = { 5'd1,	5'd4,	5'd18,	5'd9};
		rom[ 2607 ] = { 5'd15,	5'd12,	5'd9,	5'd6};
		rom[ 2608 ] = { 5'd3,	5'd9,	5'd18,	5'd6};
		rom[ 2609 ] = { 5'd18,	5'd5,	5'd6,	5'd9};
		rom[ 2610 ] = { 5'd0,	5'd5,	5'd6,	5'd9};
		rom[ 2611 ] = { 5'd4,	5'd7,	5'd18,	5'd4};
		rom[ 2612 ] = { 5'd2,	5'd1,	5'd12,	5'd20};
		rom[ 2613 ] = { 5'd17,	5'd0,	5'd6,	5'd23};
		rom[ 2614 ] = { 5'd1,	5'd6,	5'd2,	5'd18};
		rom[ 2615 ] = { 5'd8,	5'd8,	5'd10,	5'd6};
		rom[ 2616 ] = { 5'd0,	5'd6,	5'd20,	5'd6};
		rom[ 2617 ] = { 5'd11,	5'd12,	5'd12,	5'd5};
		rom[ 2618 ] = { 5'd0,	5'd4,	5'd3,	5'd19};
		rom[ 2619 ] = { 5'd19,	5'd1,	5'd3,	5'd18};
		rom[ 2620 ] = { 5'd2,	5'd1,	5'd3,	5'd18};
		rom[ 2621 ] = { 5'd3,	5'd10,	5'd18,	5'd3};
		rom[ 2622 ] = { 5'd4,	5'd4,	5'd10,	5'd9};
		rom[ 2623 ] = { 5'd7,	5'd13,	5'd14,	5'd7};
		rom[ 2624 ] = { 5'd3,	5'd13,	5'd14,	5'd7};
		rom[ 2625 ] = { 5'd8,	5'd15,	5'd9,	5'd6};
		rom[ 2626 ] = { 5'd4,	5'd14,	5'd8,	5'd10};
		rom[ 2627 ] = { 5'd10,	5'd14,	5'd4,	5'd10};
		rom[ 2628 ] = { 5'd3,	5'd8,	5'd5,	5'd16};
		rom[ 2629 ] = { 5'd15,	5'd10,	5'd9,	5'd6};
		rom[ 2630 ] = { 5'd0,	5'd10,	5'd9,	5'd6};
		rom[ 2631 ] = { 5'd6,	5'd7,	5'd12,	5'd9};
		rom[ 2632 ] = { 5'd9,	5'd10,	5'd5,	5'd8};
		rom[ 2633 ] = { 5'd12,	5'd1,	5'd3,	5'd12};
		rom[ 2634 ] = { 5'd8,	5'd15,	5'd6,	5'd9};
		rom[ 2635 ] = { 5'd16,	5'd6,	5'd7,	5'd6};
		rom[ 2636 ] = { 5'd8,	5'd1,	5'd4,	5'd22};
		rom[ 2637 ] = { 5'd6,	5'd6,	5'd14,	5'd3};
		rom[ 2638 ] = { 5'd0,	5'd18,	5'd19,	5'd3};
		rom[ 2639 ] = { 5'd17,	5'd0,	5'd6,	5'd24};
		rom[ 2640 ] = { 5'd0,	5'd13,	5'd15,	5'd6};
		rom[ 2641 ] = { 5'd9,	5'd6,	5'd10,	5'd14};
		rom[ 2642 ] = { 5'd1,	5'd6,	5'd8,	5'd10};
		rom[ 2643 ] = { 5'd7,	5'd6,	5'd12,	5'd5};
		rom[ 2644 ] = { 5'd7,	5'd7,	5'd9,	5'd6};
		rom[ 2645 ] = { 5'd7,	5'd8,	5'd14,	5'd14};
		rom[ 2646 ] = { 5'd3,	5'd8,	5'd14,	5'd14};
		rom[ 2647 ] = { 5'd9,	5'd8,	5'd13,	5'd4};
		rom[ 2648 ] = { 5'd3,	5'd2,	5'd6,	5'd12};
		rom[ 2649 ] = { 5'd6,	5'd10,	5'd17,	5'd6};
		rom[ 2650 ] = { 5'd1,	5'd10,	5'd17,	5'd6};
		rom[ 2651 ] = { 5'd16,	5'd7,	5'd8,	5'd9};
		rom[ 2652 ] = { 5'd0,	5'd7,	5'd8,	5'd9};
		rom[ 2653 ] = { 5'd0,	5'd9,	5'd24,	5'd10};
		rom[ 2654 ] = { 5'd3,	5'd2,	5'd15,	5'd8};
		rom[ 2655 ] = { 5'd4,	5'd2,	5'd18,	5'd8};
		rom[ 2656 ] = { 5'd0,	5'd1,	5'd18,	5'd4};
		rom[ 2657 ] = { 5'd20,	5'd2,	5'd3,	5'd18};
		rom[ 2658 ] = { 5'd1,	5'd3,	5'd3,	5'd19};
		rom[ 2659 ] = { 5'd18,	5'd8,	5'd6,	5'd16};
		rom[ 2660 ] = { 5'd0,	5'd8,	5'd6,	5'd16};
		rom[ 2661 ] = { 5'd8,	5'd18,	5'd11,	5'd6};
		rom[ 2662 ] = { 5'd4,	5'd6,	5'd12,	5'd5};
		rom[ 2663 ] = { 5'd7,	5'd6,	5'd12,	5'd5};
		rom[ 2664 ] = { 5'd6,	5'd3,	5'd9,	5'd6};
		rom[ 2665 ] = { 5'd7,	5'd6,	5'd12,	5'd5};
		rom[ 2666 ] = { 5'd9,	5'd8,	5'd6,	5'd7};
		rom[ 2667 ] = { 5'd8,	5'd2,	5'd9,	5'd6};
		rom[ 2668 ] = { 5'd8,	5'd14,	5'd6,	5'd9};
		rom[ 2669 ] = { 5'd8,	5'd2,	5'd9,	5'd6};
		rom[ 2670 ] = { 5'd4,	5'd3,	5'd16,	5'd20};
		rom[ 2671 ] = { 5'd7,	5'd6,	5'd10,	5'd12};
		rom[ 2672 ] = { 5'd0,	5'd2,	5'd7,	5'd12};
		rom[ 2673 ] = { 5'd12,	5'd17,	5'd11,	5'd6};
		rom[ 2674 ] = { 5'd4,	5'd7,	5'd12,	5'd8};
		rom[ 2675 ] = { 5'd8,	5'd11,	5'd8,	5'd10};
		rom[ 2676 ] = { 5'd9,	5'd1,	5'd4,	5'd9};
		rom[ 2677 ] = { 5'd14,	5'd0,	5'd3,	5'd22};
		rom[ 2678 ] = { 5'd7,	5'd0,	5'd3,	5'd22};
		rom[ 2679 ] = { 5'd4,	5'd7,	5'd18,	5'd4};
		rom[ 2680 ] = { 5'd10,	5'd2,	5'd4,	5'd15};
		rom[ 2681 ] = { 5'd12,	5'd1,	5'd3,	5'd12};
		rom[ 2682 ] = { 5'd0,	5'd0,	5'd18,	5'd13};
		rom[ 2683 ] = { 5'd16,	5'd0,	5'd3,	5'd24};
		rom[ 2684 ] = { 5'd5,	5'd0,	5'd3,	5'd24};
		rom[ 2685 ] = { 5'd10,	5'd15,	5'd5,	5'd8};
		rom[ 2686 ] = { 5'd2,	5'd18,	5'd18,	5'd2};
		rom[ 2687 ] = { 5'd2,	5'd8,	5'd20,	5'd3};
		rom[ 2688 ] = { 5'd7,	5'd6,	5'd9,	5'd6};
		rom[ 2689 ] = { 5'd3,	5'd2,	5'd19,	5'd10};
		rom[ 2690 ] = { 5'd2,	5'd7,	5'd19,	5'd3};
		rom[ 2691 ] = { 5'd15,	5'd6,	5'd9,	5'd4};
		rom[ 2692 ] = { 5'd2,	5'd2,	5'd18,	5'd8};
		rom[ 2693 ] = { 5'd10,	5'd9,	5'd14,	5'd4};
		rom[ 2694 ] = { 5'd4,	5'd4,	5'd6,	5'd16};
		rom[ 2695 ] = { 5'd15,	5'd8,	5'd9,	5'd16};
		rom[ 2696 ] = { 5'd0,	5'd8,	5'd9,	5'd16};
		rom[ 2697 ] = { 5'd18,	5'd0,	5'd6,	5'd14};
		rom[ 2698 ] = { 5'd0,	5'd0,	5'd6,	5'd14};
		rom[ 2699 ] = { 5'd15,	5'd0,	5'd6,	5'd22};
		rom[ 2700 ] = { 5'd3,	5'd0,	5'd6,	5'd22};
		rom[ 2701 ] = { 5'd12,	5'd2,	5'd12,	5'd20};
		rom[ 2702 ] = { 5'd0,	5'd2,	5'd12,	5'd20};
		rom[ 2703 ] = { 5'd11,	5'd6,	5'd4,	5'd9};
		rom[ 2704 ] = { 5'd9,	5'd0,	5'd6,	5'd16};
		rom[ 2705 ] = { 5'd12,	5'd1,	5'd3,	5'd12};
		rom[ 2706 ] = { 5'd3,	5'd4,	5'd18,	5'd6};
		rom[ 2707 ] = { 5'd5,	5'd5,	5'd16,	5'd8};
		rom[ 2708 ] = { 5'd0,	5'd13,	5'd10,	5'd6};
		rom[ 2709 ] = { 5'd8,	5'd14,	5'd9,	5'd6};
		rom[ 2710 ] = { 5'd6,	5'd2,	5'd9,	5'd6};
		rom[ 2711 ] = { 5'd14,	5'd1,	5'd10,	5'd8};
		rom[ 2712 ] = { 5'd9,	5'd1,	5'd3,	5'd12};
		rom[ 2713 ] = { 5'd6,	5'd4,	5'd12,	5'd9};
		rom[ 2714 ] = { 5'd6,	5'd5,	5'd12,	5'd6};
		rom[ 2715 ] = { 5'd1,	5'd1,	5'd8,	5'd5};
		rom[ 2716 ] = { 5'd12,	5'd12,	5'd6,	5'd8};
		rom[ 2717 ] = { 5'd3,	5'd12,	5'd12,	5'd6};
		rom[ 2718 ] = { 5'd9,	5'd18,	5'd12,	5'd6};
		rom[ 2719 ] = { 5'd4,	5'd13,	5'd6,	5'd6};
		rom[ 2720 ] = { 5'd11,	5'd3,	5'd7,	5'd18};
		rom[ 2721 ] = { 5'd3,	5'd9,	5'd18,	5'd3};
		rom[ 2722 ] = { 5'd5,	5'd3,	5'd19,	5'd2};
		rom[ 2723 ] = { 5'd4,	5'd2,	5'd12,	5'd6};
		rom[ 2724 ] = { 5'd9,	5'd6,	5'd6,	5'd9};
		rom[ 2725 ] = { 5'd8,	5'd6,	5'd6,	5'd9};
		rom[ 2726 ] = { 5'd16,	5'd9,	5'd5,	5'd15};
		rom[ 2727 ] = { 5'd3,	5'd9,	5'd5,	5'd15};
		rom[ 2728 ] = { 5'd6,	5'd6,	5'd14,	5'd6};
		rom[ 2729 ] = { 5'd8,	5'd6,	5'd3,	5'd14};
		rom[ 2730 ] = { 5'd0,	5'd16,	5'd24,	5'd5};
		rom[ 2731 ] = { 5'd0,	5'd20,	5'd20,	5'd3};
		rom[ 2732 ] = { 5'd5,	5'd10,	5'd18,	5'd2};
		rom[ 2733 ] = { 5'd0,	5'd6,	5'd6,	5'd10};
		rom[ 2734 ] = { 5'd2,	5'd1,	5'd20,	5'd3};
		rom[ 2735 ] = { 5'd9,	5'd13,	5'd6,	5'd11};
		rom[ 2736 ] = { 5'd9,	5'd15,	5'd6,	5'd8};
		rom[ 2737 ] = { 5'd9,	5'd12,	5'd6,	5'd9};
		rom[ 2738 ] = { 5'd5,	5'd11,	5'd18,	5'd2};
		rom[ 2739 ] = { 5'd2,	5'd6,	5'd15,	5'd6};
		rom[ 2740 ] = { 5'd6,	5'd0,	5'd18,	5'd3};
		rom[ 2741 ] = { 5'd5,	5'd0,	5'd3,	5'd18};
		rom[ 2742 ] = { 5'd18,	5'd3,	5'd6,	5'd10};
		rom[ 2743 ] = { 5'd0,	5'd3,	5'd6,	5'd10};
		rom[ 2744 ] = { 5'd10,	5'd5,	5'd8,	5'd9};
		rom[ 2745 ] = { 5'd6,	5'd5,	5'd8,	5'd9};
		rom[ 2746 ] = { 5'd3,	5'd2,	5'd20,	5'd3};
		rom[ 2747 ] = { 5'd5,	5'd2,	5'd13,	5'd4};
		rom[ 2748 ] = { 5'd17,	5'd0,	5'd7,	5'd14};
		rom[ 2749 ] = { 5'd0,	5'd0,	5'd7,	5'd14};
		rom[ 2750 ] = { 5'd9,	5'd11,	5'd10,	5'd6};
		rom[ 2751 ] = { 5'd5,	5'd11,	5'd10,	5'd6};
		rom[ 2752 ] = { 5'd11,	5'd6,	5'd3,	5'd18};
		rom[ 2753 ] = { 5'd0,	5'd16,	5'd18,	5'd3};
		rom[ 2754 ] = { 5'd6,	5'd16,	5'd18,	5'd3};
		rom[ 2755 ] = { 5'd4,	5'd6,	5'd9,	5'd10};
		rom[ 2756 ] = { 5'd9,	5'd7,	5'd15,	5'd4};
		rom[ 2757 ] = { 5'd5,	5'd6,	5'd12,	5'd6};
		rom[ 2758 ] = { 5'd6,	5'd1,	5'd12,	5'd9};
		rom[ 2759 ] = { 5'd7,	5'd9,	5'd6,	5'd12};
		rom[ 2760 ] = { 5'd11,	5'd5,	5'd13,	5'd6};
		rom[ 2761 ] = { 5'd1,	5'd11,	5'd22,	5'd13};
		rom[ 2762 ] = { 5'd18,	5'd8,	5'd6,	5'd6};
		rom[ 2763 ] = { 5'd0,	5'd8,	5'd6,	5'd6};
		rom[ 2764 ] = { 5'd0,	5'd6,	5'd24,	5'd3};
		rom[ 2765 ] = { 5'd0,	5'd5,	5'd10,	5'd6};
		rom[ 2766 ] = { 5'd6,	5'd7,	5'd18,	5'd3};
		rom[ 2767 ] = { 5'd0,	5'd0,	5'd10,	5'd6};
		rom[ 2768 ] = { 5'd19,	5'd0,	5'd3,	5'd19};
		rom[ 2769 ] = { 5'd4,	5'd6,	5'd12,	5'd16};
		rom[ 2770 ] = { 5'd19,	5'd6,	5'd4,	5'd18};
		rom[ 2771 ] = { 5'd1,	5'd6,	5'd4,	5'd18};
		rom[ 2772 ] = { 5'd3,	5'd21,	5'd18,	5'd3};
		rom[ 2773 ] = { 5'd0,	5'd19,	5'd9,	5'd4};
		rom[ 2774 ] = { 5'd12,	5'd18,	5'd12,	5'd6};
		rom[ 2775 ] = { 5'd7,	5'd18,	5'd9,	5'd4};
		rom[ 2776 ] = { 5'd12,	5'd16,	5'd10,	5'd8};
		rom[ 2777 ] = { 5'd2,	5'd16,	5'd10,	5'd8};
		rom[ 2778 ] = { 5'd14,	5'd0,	5'd10,	5'd12};
		rom[ 2779 ] = { 5'd0,	5'd0,	5'd10,	5'd12};
		rom[ 2780 ] = { 5'd15,	5'd14,	5'd9,	5'd6};
		rom[ 2781 ] = { 5'd0,	5'd14,	5'd9,	5'd6};
		rom[ 2782 ] = { 5'd14,	5'd14,	5'd10,	5'd6};
		rom[ 2783 ] = { 5'd0,	5'd14,	5'd10,	5'd6};
		rom[ 2784 ] = { 5'd5,	5'd18,	5'd18,	5'd2};
		rom[ 2785 ] = { 5'd0,	5'd18,	5'd18,	5'd3};
		rom[ 2786 ] = { 5'd3,	5'd5,	5'd18,	5'd12};
		rom[ 2787 ] = { 5'd5,	5'd3,	5'd7,	5'd9};
		rom[ 2788 ] = { 5'd4,	5'd0,	5'd19,	5'd15};
		rom[ 2789 ] = { 5'd3,	5'd0,	5'd16,	5'd4};
		rom[ 2790 ] = { 5'd4,	5'd12,	5'd16,	5'd12};
		rom[ 2791 ] = { 5'd4,	5'd3,	5'd12,	5'd15};
		rom[ 2792 ] = { 5'd16,	5'd4,	5'd2,	5'd19};
		rom[ 2793 ] = { 5'd6,	5'd4,	5'd2,	5'd19};
		rom[ 2794 ] = { 5'd13,	5'd14,	5'd8,	5'd10};
		rom[ 2795 ] = { 5'd3,	5'd14,	5'd8,	5'd10};
		rom[ 2796 ] = { 5'd12,	5'd6,	5'd3,	5'd18};
		rom[ 2797 ] = { 5'd5,	5'd11,	5'd12,	5'd6};
		rom[ 2798 ] = { 5'd10,	5'd5,	5'd8,	5'd10};
		rom[ 2799 ] = { 5'd6,	5'd4,	5'd12,	5'd10};
		rom[ 2800 ] = { 5'd6,	5'd8,	5'd18,	5'd10};
		rom[ 2801 ] = { 5'd0,	5'd8,	5'd18,	5'd10};
		rom[ 2802 ] = { 5'd12,	5'd6,	5'd3,	5'd18};
		rom[ 2803 ] = { 5'd0,	5'd14,	5'd18,	5'd3};
		rom[ 2804 ] = { 5'd12,	5'd6,	5'd3,	5'd18};
		rom[ 2805 ] = { 5'd9,	5'd6,	5'd3,	5'd18};
		rom[ 2806 ] = { 5'd6,	5'd14,	5'd18,	5'd3};
		rom[ 2807 ] = { 5'd0,	5'd5,	5'd18,	5'd3};
		rom[ 2808 ] = { 5'd2,	5'd5,	5'd22,	5'd3};
		rom[ 2809 ] = { 5'd0,	5'd0,	5'd21,	5'd10};
		rom[ 2810 ] = { 5'd6,	5'd3,	5'd18,	5'd17};
		rom[ 2811 ] = { 5'd0,	5'd3,	5'd18,	5'd17};
		rom[ 2812 ] = { 5'd0,	5'd12,	5'd24,	5'd11};
		rom[ 2813 ] = { 5'd4,	5'd10,	5'd16,	5'd6};
		rom[ 2814 ] = { 5'd12,	5'd8,	5'd6,	5'd8};
		rom[ 2815 ] = { 5'd6,	5'd14,	5'd8,	5'd7};
		rom[ 2816 ] = { 5'd15,	5'd10,	5'd6,	5'd14};
		rom[ 2817 ] = { 5'd3,	5'd10,	5'd6,	5'd14};
		rom[ 2818 ] = { 5'd6,	5'd12,	5'd18,	5'd2};
		rom[ 2819 ] = { 5'd5,	5'd8,	5'd10,	5'd6};
		rom[ 2820 ] = { 5'd12,	5'd11,	5'd9,	5'd4};
		rom[ 2821 ] = { 5'd0,	5'd11,	5'd9,	5'd6};
		rom[ 2822 ] = { 5'd11,	5'd2,	5'd3,	5'd18};
		rom[ 2823 ] = { 5'd10,	5'd2,	5'd3,	5'd18};
		rom[ 2824 ] = { 5'd9,	5'd12,	5'd6,	5'd10};
		rom[ 2825 ] = { 5'd1,	5'd10,	5'd6,	5'd9};
		rom[ 2826 ] = { 5'd6,	5'd9,	5'd16,	5'd6};
		rom[ 2827 ] = { 5'd1,	5'd8,	5'd9,	5'd6};
		rom[ 2828 ] = { 5'd7,	5'd7,	5'd16,	5'd6};
		rom[ 2829 ] = { 5'd0,	5'd0,	5'd18,	5'd3};
		rom[ 2830 ] = { 5'd10,	5'd0,	5'd6,	5'd9};
		rom[ 2831 ] = { 5'd9,	5'd5,	5'd6,	5'd6};
		rom[ 2832 ] = { 5'd10,	5'd6,	5'd4,	5'd18};
		rom[ 2833 ] = { 5'd8,	5'd0,	5'd6,	5'd9};
		rom[ 2834 ] = { 5'd9,	5'd1,	5'd6,	5'd9};
		rom[ 2835 ] = { 5'd1,	5'd0,	5'd18,	5'd9};
		rom[ 2836 ] = { 5'd0,	5'd3,	5'd24,	5'd3};
		rom[ 2837 ] = { 5'd6,	5'd14,	5'd9,	5'd4};
		rom[ 2838 ] = { 5'd8,	5'd9,	5'd8,	5'd10};
		rom[ 2839 ] = { 5'd5,	5'd2,	5'd13,	5'd9};
		rom[ 2840 ] = { 5'd4,	5'd4,	5'd16,	5'd9};
		rom[ 2841 ] = { 5'd4,	5'd4,	5'd14,	5'd9};
		rom[ 2842 ] = { 5'd8,	5'd5,	5'd9,	5'd6};
		rom[ 2843 ] = { 5'd1,	5'd7,	5'd16,	5'd6};
		rom[ 2844 ] = { 5'd10,	5'd5,	5'd13,	5'd9};
		rom[ 2845 ] = { 5'd1,	5'd5,	5'd13,	5'd9};
		rom[ 2846 ] = { 5'd0,	5'd4,	5'd24,	5'd6};
		rom[ 2847 ] = { 5'd1,	5'd14,	5'd10,	5'd9};
		rom[ 2848 ] = { 5'd5,	5'd17,	5'd18,	5'd3};
		rom[ 2849 ] = { 5'd0,	5'd16,	5'd18,	5'd3};
		rom[ 2850 ] = { 5'd9,	5'd17,	5'd9,	5'd6};
		rom[ 2851 ] = { 5'd1,	5'd20,	5'd22,	5'd4};
		rom[ 2852 ] = { 5'd8,	5'd14,	5'd8,	5'd6};
		rom[ 2853 ] = { 5'd8,	5'd6,	5'd8,	5'd15};
		rom[ 2854 ] = { 5'd5,	5'd4,	5'd18,	5'd3};
		rom[ 2855 ] = { 5'd9,	5'd3,	5'd5,	5'd10};
		rom[ 2856 ] = { 5'd6,	5'd8,	5'd12,	5'd3};
		rom[ 2857 ] = { 5'd2,	5'd6,	5'd18,	5'd6};
		rom[ 2858 ] = { 5'd10,	5'd6,	5'd4,	5'd18};
		rom[ 2859 ] = { 5'd7,	5'd5,	5'd6,	5'd6};
		rom[ 2860 ] = { 5'd14,	5'd5,	5'd2,	5'd18};
		rom[ 2861 ] = { 5'd8,	5'd5,	5'd2,	5'd18};
		rom[ 2862 ] = { 5'd9,	5'd2,	5'd10,	5'd6};
		rom[ 2863 ] = { 5'd3,	5'd1,	5'd18,	5'd12};
		rom[ 2864 ] = { 5'd5,	5'd2,	5'd17,	5'd22};
		rom[ 2865 ] = { 5'd4,	5'd0,	5'd12,	5'd6};
		rom[ 2866 ] = { 5'd6,	5'd9,	5'd16,	5'd6};
		rom[ 2867 ] = { 5'd9,	5'd0,	5'd5,	5'd18};
		rom[ 2868 ] = { 5'd12,	5'd0,	5'd6,	5'd9};
		rom[ 2869 ] = { 5'd6,	5'd0,	5'd6,	5'd9};
		rom[ 2870 ] = { 5'd9,	5'd1,	5'd6,	5'd12};
		rom[ 2871 ] = { 5'd5,	5'd9,	5'd13,	5'd4};
		rom[ 2872 ] = { 5'd5,	5'd8,	5'd19,	5'd3};
		rom[ 2873 ] = { 5'd9,	5'd9,	5'd6,	5'd8};
		rom[ 2874 ] = { 5'd11,	5'd9,	5'd4,	5'd15};
		rom[ 2875 ] = { 5'd2,	5'd0,	5'd6,	5'd14};
		rom[ 2876 ] = { 5'd15,	5'd1,	5'd6,	5'd14};
		rom[ 2877 ] = { 5'd3,	5'd1,	5'd6,	5'd14};
		rom[ 2878 ] = { 5'd3,	5'd20,	5'd18,	5'd4};
		rom[ 2879 ] = { 5'd5,	5'd0,	5'd4,	5'd20};
		rom[ 2880 ] = { 5'd16,	5'd8,	5'd8,	5'd12};
		rom[ 2881 ] = { 5'd0,	5'd8,	5'd8,	5'd12};
		rom[ 2882 ] = { 5'd13,	5'd13,	5'd10,	5'd8};
		rom[ 2883 ] = { 5'd1,	5'd13,	5'd10,	5'd8};
		rom[ 2884 ] = { 5'd15,	5'd8,	5'd4,	5'd15};
		rom[ 2885 ] = { 5'd5,	5'd8,	5'd4,	5'd15};
		rom[ 2886 ] = { 5'd6,	5'd11,	5'd16,	5'd12};
		rom[ 2887 ] = { 5'd2,	5'd11,	5'd16,	5'd12};
		rom[ 2888 ] = { 5'd14,	5'd12,	5'd7,	5'd9};
		rom[ 2889 ] = { 5'd10,	5'd1,	5'd3,	5'd21};
		rom[ 2890 ] = { 5'd13,	5'd11,	5'd9,	5'd4};
		rom[ 2891 ] = { 5'd3,	5'd10,	5'd17,	5'd9};
		rom[ 2892 ] = { 5'd13,	5'd8,	5'd8,	5'd15};
		rom[ 2893 ] = { 5'd3,	5'd8,	5'd8,	5'd15};
		rom[ 2894 ] = { 5'd11,	5'd14,	5'd10,	5'd8};
		rom[ 2895 ] = { 5'd0,	5'd18,	5'd22,	5'd6};
		rom[ 2896 ] = { 5'd0,	5'd16,	5'd24,	5'd4};
		rom[ 2897 ] = { 5'd6,	5'd20,	5'd12,	5'd3};
		rom[ 2898 ] = { 5'd18,	5'd12,	5'd6,	5'd12};
		rom[ 2899 ] = { 5'd0,	5'd12,	5'd6,	5'd12};
		rom[ 2900 ] = { 5'd15,	5'd17,	5'd9,	5'd6};
		rom[ 2901 ] = { 5'd1,	5'd6,	5'd22,	5'd10};
		rom[ 2902 ] = { 5'd15,	5'd17,	5'd9,	5'd6};
		rom[ 2903 ] = { 5'd0,	5'd18,	5'd18,	5'd2};
		rom[ 2904 ] = { 5'd3,	5'd15,	5'd19,	5'd3};
		rom[ 2905 ] = { 5'd0,	5'd13,	5'd18,	5'd3};
		rom[ 2906 ] = { 5'd15,	5'd17,	5'd9,	5'd6};
		rom[ 2907 ] = { 5'd0,	5'd17,	5'd9,	5'd6};
		rom[ 2908 ] = { 5'd12,	5'd17,	5'd9,	5'd6};
		rom[ 2909 ] = { 5'd3,	5'd17,	5'd9,	5'd6};
		rom[ 2910 ] = { 5'd16,	5'd2,	5'd3,	5'd20};
		rom[ 2911 ] = { 5'd0,	5'd13,	5'd24,	5'd8};
		rom[ 2912 ] = { 5'd9,	5'd1,	5'd6,	5'd22};

	end
endmodule


module rect1_rom(
	input 				clk,
	input		[11:0]	addr,
	output reg	[19:0]	q    // x y w h 5bit*4
	);
	reg					[19:0]	rom [4095:0];
	always @(posedge clk) q <= rom[addr];
	initial begin
		rom[ 0    ] = { 5'd6,	5'd7,	5'd12,	5'd3};
		rom[ 1    ] = { 5'd10,	5'd4,	5'd4,	5'd7};
		rom[ 2    ] = { 5'd3,	5'd12,	5'd18,	5'd3};
		rom[ 3    ] = { 5'd8,	5'd20,	5'd9,	5'd2};
		rom[ 4    ] = { 5'd5,	5'd5,	5'd2,	5'd19};
		rom[ 5    ] = { 5'd6,	5'd13,	5'd12,	5'd8};
		rom[ 6    ] = { 5'd5,	5'd11,	5'd12,	5'd3};
		rom[ 7    ] = { 5'd11,	5'd19,	5'd4,	5'd5};
		rom[ 8    ] = { 5'd4,	5'd3,	5'd7,	5'd3};
		rom[ 9    ] = { 5'd6,	5'd8,	5'd12,	5'd2};
		rom[ 10   ] = { 5'd10,	5'd4,	5'd4,	5'd7};
		rom[ 11   ] = { 5'd1,	5'd12,	5'd19,	5'd4};
		rom[ 12   ] = { 5'd8,	5'd2,	5'd8,	5'd3};
		rom[ 13   ] = { 5'd9,	5'd14,	5'd6,	5'd5};
		rom[ 14   ] = { 5'd5,	5'd11,	5'd14,	5'd5};
		rom[ 15   ] = { 5'd5,	5'd3,	5'd14,	5'd3};
		rom[ 16   ] = { 5'd16,	5'd11,	5'd3,	5'd6};
		rom[ 17   ] = { 5'd9,	5'd5,	5'd2,	5'd10};
		rom[ 18   ] = { 5'd12,	5'd8,	5'd2,	5'd10};
		rom[ 19   ] = { 5'd4,	5'd5,	5'd2,	5'd9};
		rom[ 20   ] = { 5'd20,	5'd0,	5'd2,	5'd11};
		rom[ 21   ] = { 5'd8,	5'd6,	5'd8,	5'd13};
		rom[ 22   ] = { 5'd11,	5'd6,	5'd2,	5'd9};
		rom[ 23   ] = { 5'd7,	5'd20,	5'd10,	5'd2};
		rom[ 24   ] = { 5'd5,	5'd13,	5'd14,	5'd6};
		rom[ 25   ] = { 5'd8,	5'd3,	5'd8,	5'd3};
		rom[ 26   ] = { 5'd5,	5'd11,	5'd15,	5'd3};
		rom[ 27   ] = { 5'd9,	5'd13,	5'd5,	5'd7};
		rom[ 28   ] = { 5'd11,	5'd5,	5'd2,	5'd10};
		rom[ 29   ] = { 5'd6,	5'd12,	5'd3,	5'd6};
		rom[ 30   ] = { 5'd9,	5'd21,	5'd6,	5'd3};
		rom[ 31   ] = { 5'd5,	5'd8,	5'd13,	5'd2};
		rom[ 32   ] = { 5'd18,	5'd1,	5'd3,	5'd15};
		rom[ 33   ] = { 5'd4,	5'd1,	5'd3,	5'd15};
		rom[ 34   ] = { 5'd8,	5'd8,	5'd8,	5'd15};
		rom[ 35   ] = { 5'd5,	5'd6,	5'd7,	5'd6};
		rom[ 36   ] = { 5'd2,	5'd16,	5'd21,	5'd4};
		rom[ 37   ] = { 5'd10,	5'd1,	5'd2,	5'd10};
		rom[ 38   ] = { 5'd2,	5'd13,	5'd10,	5'd10};
		rom[ 39   ] = { 5'd2,	5'd1,	5'd2,	5'd13};
		rom[ 40   ] = { 5'd20,	5'd2,	5'd2,	5'd13};
		rom[ 41   ] = { 5'd11,	5'd5,	5'd11,	5'd19};
		rom[ 42   ] = { 5'd20,	5'd4,	5'd2,	5'd9};
		rom[ 43   ] = { 5'd2,	5'd3,	5'd2,	5'd11};
		rom[ 44   ] = { 5'd12,	5'd1,	5'd2,	5'd9};
		rom[ 45   ] = { 5'd0,	5'd7,	5'd19,	5'd1};
		rom[ 46   ] = { 5'd12,	5'd1,	5'd2,	5'd9};
		rom[ 47   ] = { 5'd10,	5'd1,	5'd2,	5'd9};
		rom[ 48   ] = { 5'd12,	5'd5,	5'd7,	5'd7};
		rom[ 49   ] = { 5'd1,	5'd11,	5'd18,	5'd1};
		rom[ 50   ] = { 5'd17,	5'd13,	5'd2,	5'd11};
		rom[ 51   ] = { 5'd0,	5'd7,	5'd6,	5'd3};
		rom[ 52   ] = { 5'd6,	5'd7,	5'd12,	5'd3};
		rom[ 53   ] = { 5'd10,	5'd5,	5'd4,	5'd6};
		rom[ 54   ] = { 5'd8,	5'd1,	5'd8,	5'd5};
		rom[ 55   ] = { 5'd4,	5'd12,	5'd18,	5'd2};
		rom[ 56   ] = { 5'd2,	5'd17,	5'd6,	5'd3};
		rom[ 57   ] = { 5'd19,	5'd3,	5'd2,	5'd13};
		rom[ 58   ] = { 5'd3,	5'd3,	5'd2,	5'd13};
		rom[ 59   ] = { 5'd8,	5'd1,	5'd8,	5'd23};
		rom[ 60   ] = { 5'd1,	5'd11,	5'd8,	5'd4};
		rom[ 61   ] = { 5'd14,	5'd14,	5'd3,	5'd7};
		rom[ 62   ] = { 5'd3,	5'd12,	5'd8,	5'd3};
		rom[ 63   ] = { 5'd6,	5'd8,	5'd12,	5'd2};
		rom[ 64   ] = { 5'd8,	5'd13,	5'd6,	5'd6};
		rom[ 65   ] = { 5'd15,	5'd17,	5'd9,	5'd2};
		rom[ 66   ] = { 5'd1,	5'd18,	5'd18,	5'd1};
		rom[ 67   ] = { 5'd4,	5'd10,	5'd16,	5'd6};
		rom[ 68   ] = { 5'd2,	5'd1,	5'd2,	5'd20};
		rom[ 69   ] = { 5'd3,	5'd1,	5'd18,	5'd1};
		rom[ 70   ] = { 5'd1,	5'd5,	5'd10,	5'd7};
		rom[ 71   ] = { 5'd5,	5'd12,	5'd14,	5'd4};
		rom[ 72   ] = { 5'd3,	5'd17,	5'd7,	5'd3};
		rom[ 73   ] = { 5'd14,	5'd17,	5'd9,	5'd2};
		rom[ 74   ] = { 5'd1,	5'd17,	5'd9,	5'd2};
		rom[ 75   ] = { 5'd15,	5'd6,	5'd4,	5'd5};
		rom[ 76   ] = { 5'd5,	5'd5,	5'd7,	5'd7};
		rom[ 77   ] = { 5'd10,	5'd0,	5'd4,	5'd5};
		rom[ 78   ] = { 5'd9,	5'd3,	5'd6,	5'd3};
		rom[ 79   ] = { 5'd11,	5'd6,	5'd2,	5'd9};
		rom[ 80   ] = { 5'd9,	5'd0,	5'd2,	5'd9};
		rom[ 81   ] = { 5'd12,	5'd6,	5'd2,	5'd9};
		rom[ 82   ] = { 5'd10,	5'd6,	5'd2,	5'd9};
		rom[ 83   ] = { 5'd9,	5'd8,	5'd6,	5'd4};
		rom[ 84   ] = { 5'd6,	5'd3,	5'd12,	5'd3};
		rom[ 85   ] = { 5'd8,	5'd0,	5'd8,	5'd6};
		rom[ 86   ] = { 5'd4,	5'd11,	5'd16,	5'd4};
		rom[ 87   ] = { 5'd11,	5'd6,	5'd3,	5'd6};
		rom[ 88   ] = { 5'd8,	5'd20,	5'd8,	5'd3};
		rom[ 89   ] = { 5'd11,	5'd6,	5'd2,	5'd9};
		rom[ 90   ] = { 5'd9,	5'd13,	5'd5,	5'd4};
		rom[ 91   ] = { 5'd11,	5'd6,	5'd2,	5'd9};
		rom[ 92   ] = { 5'd11,	5'd6,	5'd2,	5'd9};
		rom[ 93   ] = { 5'd9,	5'd18,	5'd6,	5'd6};
		rom[ 94   ] = { 5'd1,	5'd23,	5'd18,	5'd1};
		rom[ 95   ] = { 5'd10,	5'd12,	5'd4,	5'd5};
		rom[ 96   ] = { 5'd6,	5'd12,	5'd8,	5'd5};
		rom[ 97   ] = { 5'd7,	5'd8,	5'd10,	5'd2};
		rom[ 98   ] = { 5'd0,	5'd16,	5'd10,	5'd2};
		rom[ 99   ] = { 5'd6,	5'd19,	5'd18,	5'd1};
		rom[ 100  ] = { 5'd1,	5'd2,	5'd22,	5'd1};
		rom[ 101  ] = { 5'd6,	5'd17,	5'd18,	5'd1};
		rom[ 102  ] = { 5'd5,	5'd4,	5'd3,	5'd15};
		rom[ 103  ] = { 5'd20,	5'd4,	5'd2,	5'd10};
		rom[ 104  ] = { 5'd2,	5'd4,	5'd2,	5'd10};
		rom[ 105  ] = { 5'd12,	5'd16,	5'd10,	5'd3};
		rom[ 106  ] = { 5'd4,	5'd12,	5'd4,	5'd9};
		rom[ 107  ] = { 5'd14,	5'd0,	5'd2,	5'd9};
		rom[ 108  ] = { 5'd8,	5'd10,	5'd3,	5'd6};
		rom[ 109  ] = { 5'd17,	5'd8,	5'd6,	5'd3};
		rom[ 110  ] = { 5'd0,	5'd8,	5'd6,	5'd3};
		rom[ 111  ] = { 5'd14,	5'd0,	5'd2,	5'd9};
		rom[ 112  ] = { 5'd8,	5'd0,	5'd2,	5'd9};
		rom[ 113  ] = { 5'd8,	5'd16,	5'd9,	5'd2};
		rom[ 114  ] = { 5'd0,	5'd18,	5'd9,	5'd2};
		rom[ 115  ] = { 5'd12,	5'd8,	5'd2,	5'd10};
		rom[ 116  ] = { 5'd9,	5'd19,	5'd6,	5'd3};
		rom[ 117  ] = { 5'd2,	5'd11,	5'd20,	5'd1};
		rom[ 118  ] = { 5'd2,	5'd9,	5'd9,	5'd6};
		rom[ 119  ] = { 5'd3,	5'd0,	5'd9,	5'd24};
		rom[ 120  ] = { 5'd5,	5'd6,	5'd7,	5'd5};
		rom[ 121  ] = { 5'd14,	5'd5,	5'd5,	5'd6};
		rom[ 122  ] = { 5'd4,	5'd5,	5'd6,	5'd6};
		rom[ 123  ] = { 5'd4,	5'd15,	5'd18,	5'd1};
		rom[ 124  ] = { 5'd6,	5'd17,	5'd8,	5'd4};
		rom[ 125  ] = { 5'd3,	5'd19,	5'd18,	5'd3};
		rom[ 126  ] = { 5'd3,	5'd0,	5'd3,	5'd6};
		rom[ 127  ] = { 5'd10,	5'd6,	5'd4,	5'd18};
		rom[ 128  ] = { 5'd8,	5'd1,	5'd2,	5'd14};
		rom[ 129  ] = { 5'd3,	5'd3,	5'd19,	5'd1};
		rom[ 130  ] = { 5'd12,	5'd8,	5'd11,	5'd13};
		rom[ 131  ] = { 5'd8,	5'd11,	5'd11,	5'd2};
		rom[ 132  ] = { 5'd5,	5'd12,	5'd5,	5'd10};
		rom[ 133  ] = { 5'd16,	5'd16,	5'd4,	5'd6};
		rom[ 134  ] = { 5'd4,	5'd16,	5'd4,	5'd6};
		rom[ 135  ] = { 5'd19,	5'd5,	5'd5,	5'd4};
		rom[ 136  ] = { 5'd8,	5'd2,	5'd8,	5'd4};
		rom[ 137  ] = { 5'd6,	5'd10,	5'd12,	5'd2};
		rom[ 138  ] = { 5'd10,	5'd5,	5'd3,	5'd6};
		rom[ 139  ] = { 5'd9,	5'd20,	5'd6,	5'd3};
		rom[ 140  ] = { 5'd0,	5'd12,	5'd22,	5'd5};
		rom[ 141  ] = { 5'd4,	5'd4,	5'd17,	5'd3};
		rom[ 142  ] = { 5'd9,	5'd5,	5'd2,	5'd10};
		rom[ 143  ] = { 5'd18,	5'd1,	5'd3,	5'd8};
		rom[ 144  ] = { 5'd3,	5'd1,	5'd3,	5'd7};
		rom[ 145  ] = { 5'd18,	5'd0,	5'd3,	5'd22};
		rom[ 146  ] = { 5'd3,	5'd0,	5'd3,	5'd22};
		rom[ 147  ] = { 5'd16,	5'd7,	5'd4,	5'd16};
		rom[ 148  ] = { 5'd2,	5'd12,	5'd19,	5'd2};
		rom[ 149  ] = { 5'd9,	5'd13,	5'd6,	5'd4};
		rom[ 150  ] = { 5'd2,	5'd17,	5'd17,	5'd2};
		rom[ 151  ] = { 5'd14,	5'd14,	5'd3,	5'd7};
		rom[ 152  ] = { 5'd5,	5'd6,	5'd4,	5'd5};
		rom[ 153  ] = { 5'd18,	5'd8,	5'd3,	5'd11};
		rom[ 154  ] = { 5'd3,	5'd8,	5'd3,	5'd11};
		rom[ 155  ] = { 5'd8,	5'd15,	5'd10,	5'd9};
		rom[ 156  ] = { 5'd7,	5'd14,	5'd3,	5'd7};
		rom[ 157  ] = { 5'd8,	5'd14,	5'd8,	5'd8};
		rom[ 158  ] = { 5'd10,	5'd10,	5'd9,	5'd14};
		rom[ 159  ] = { 5'd14,	5'd15,	5'd6,	5'd3};
		rom[ 160  ] = { 5'd7,	5'd0,	5'd5,	5'd8};
		rom[ 161  ] = { 5'd13,	5'd0,	5'd3,	5'd6};
		rom[ 162  ] = { 5'd12,	5'd3,	5'd8,	5'd4};
		rom[ 163  ] = { 5'd13,	5'd0,	5'd3,	5'd6};
		rom[ 164  ] = { 5'd1,	5'd1,	5'd10,	5'd2};
		rom[ 165  ] = { 5'd13,	5'd0,	5'd3,	5'd6};
		rom[ 166  ] = { 5'd8,	5'd0,	5'd3,	5'd6};
		rom[ 167  ] = { 5'd8,	5'd20,	5'd10,	5'd2};
		rom[ 168  ] = { 5'd8,	5'd3,	5'd2,	5'd9};
		rom[ 169  ] = { 5'd7,	5'd5,	5'd12,	5'd2};
		rom[ 170  ] = { 5'd0,	5'd11,	5'd18,	5'd1};
		rom[ 171  ] = { 5'd1,	5'd11,	5'd22,	5'd1};
		rom[ 172  ] = { 5'd9,	5'd11,	5'd4,	5'd8};
		rom[ 173  ] = { 5'd12,	5'd11,	5'd3,	5'd6};
		rom[ 174  ] = { 5'd9,	5'd11,	5'd3,	5'd6};
		rom[ 175  ] = { 5'd7,	5'd12,	5'd11,	5'd2};
		rom[ 176  ] = { 5'd0,	5'd13,	5'd12,	5'd2};
		rom[ 177  ] = { 5'd13,	5'd4,	5'd11,	5'd6};
		rom[ 178  ] = { 5'd12,	5'd0,	5'd10,	5'd17};
		rom[ 179  ] = { 5'd14,	5'd0,	5'd1,	5'd24};
		rom[ 180  ] = { 5'd9,	5'd0,	5'd1,	5'd24};
		rom[ 181  ] = { 5'd14,	5'd1,	5'd1,	5'd22};
		rom[ 182  ] = { 5'd9,	5'd1,	5'd1,	5'd22};
		rom[ 183  ] = { 5'd18,	5'd6,	5'd1,	5'd18};
		rom[ 184  ] = { 5'd6,	5'd16,	5'd9,	5'd2};
		rom[ 185  ] = { 5'd13,	5'd16,	5'd9,	5'd2};
		rom[ 186  ] = { 5'd3,	5'd19,	5'd18,	5'd1};
		rom[ 187  ] = { 5'd13,	5'd4,	5'd4,	5'd9};
		rom[ 188  ] = { 5'd0,	5'd18,	5'd18,	5'd1};
		rom[ 189  ] = { 5'd6,	5'd2,	5'd6,	5'd4};
		rom[ 190  ] = { 5'd6,	5'd11,	5'd14,	5'd3};
		rom[ 191  ] = { 5'd10,	5'd5,	5'd3,	5'd6};
		rom[ 192  ] = { 5'd10,	5'd13,	5'd6,	5'd8};
		rom[ 193  ] = { 5'd4,	5'd4,	5'd3,	5'd16};
		rom[ 194  ] = { 5'd5,	5'd3,	5'd18,	5'd3};
		rom[ 195  ] = { 5'd9,	5'd19,	5'd5,	5'd4};
		rom[ 196  ] = { 5'd20,	5'd0,	5'd2,	5'd9};
		rom[ 197  ] = { 5'd2,	5'd1,	5'd18,	5'd1};
		rom[ 198  ] = { 5'd5,	5'd23,	5'd19,	5'd1};
		rom[ 199  ] = { 5'd2,	5'd0,	5'd2,	5'd9};
		rom[ 200  ] = { 5'd5,	5'd12,	5'd19,	5'd6};
		rom[ 201  ] = { 5'd2,	5'd1,	5'd2,	5'd9};
		rom[ 202  ] = { 5'd13,	5'd5,	5'd7,	5'd6};
		rom[ 203  ] = { 5'd0,	5'd2,	5'd20,	5'd1};
		rom[ 204  ] = { 5'd1,	5'd3,	5'd22,	5'd1};
		rom[ 205  ] = { 5'd2,	5'd11,	5'd7,	5'd3};
		rom[ 206  ] = { 5'd13,	5'd12,	5'd11,	5'd2};
		rom[ 207  ] = { 5'd0,	5'd12,	5'd11,	5'd2};
		rom[ 208  ] = { 5'd11,	5'd7,	5'd2,	5'd11};
		rom[ 209  ] = { 5'd10,	5'd1,	5'd3,	5'd6};
		rom[ 210  ] = { 5'd11,	5'd7,	5'd4,	5'd5};
		rom[ 211  ] = { 5'd6,	5'd10,	5'd12,	5'd6};
		rom[ 212  ] = { 5'd18,	5'd6,	5'd6,	5'd5};
		rom[ 213  ] = { 5'd3,	5'd16,	5'd18,	5'd1};
		rom[ 214  ] = { 5'd18,	5'd8,	5'd6,	5'd3};
		rom[ 215  ] = { 5'd1,	5'd5,	5'd8,	5'd3};
		rom[ 216  ] = { 5'd13,	5'd0,	5'd2,	5'd9};
		rom[ 217  ] = { 5'd0,	5'd4,	5'd12,	5'd7};
		rom[ 218  ] = { 5'd13,	5'd0,	5'd2,	5'd13};
		rom[ 219  ] = { 5'd9,	5'd0,	5'd2,	5'd13};
		rom[ 220  ] = { 5'd13,	5'd6,	5'd2,	5'd9};
		rom[ 221  ] = { 5'd10,	5'd7,	5'd2,	5'd9};
		rom[ 222  ] = { 5'd13,	5'd19,	5'd9,	5'd2};
		rom[ 223  ] = { 5'd2,	5'd18,	5'd7,	5'd3};
		rom[ 224  ] = { 5'd12,	5'd18,	5'd9,	5'd2};
		rom[ 225  ] = { 5'd5,	5'd20,	5'd5,	5'd4};
		rom[ 226  ] = { 5'd14,	5'd15,	5'd5,	5'd9};
		rom[ 227  ] = { 5'd4,	5'd6,	5'd16,	5'd2};
		rom[ 228  ] = { 5'd7,	5'd8,	5'd10,	5'd2};
		rom[ 229  ] = { 5'd5,	5'd14,	5'd5,	5'd10};
		rom[ 230  ] = { 5'd12,	5'd9,	5'd5,	5'd7};
		rom[ 231  ] = { 5'd9,	5'd6,	5'd2,	5'd9};
		rom[ 232  ] = { 5'd3,	5'd7,	5'd18,	5'd1};
		rom[ 233  ] = { 5'd0,	5'd11,	5'd18,	5'd1};
		rom[ 234  ] = { 5'd12,	5'd16,	5'd9,	5'd2};
		rom[ 235  ] = { 5'd4,	5'd6,	5'd7,	5'd3};
		rom[ 236  ] = { 5'd13,	5'd0,	5'd1,	5'd18};
		rom[ 237  ] = { 5'd10,	5'd0,	5'd1,	5'd18};
		rom[ 238  ] = { 5'd10,	5'd7,	5'd5,	5'd10};
		rom[ 239  ] = { 5'd8,	5'd20,	5'd7,	5'd4};
		rom[ 240  ] = { 5'd10,	5'd14,	5'd5,	5'd9};
		rom[ 241  ] = { 5'd0,	5'd2,	5'd12,	5'd3};
		rom[ 242  ] = { 5'd12,	5'd1,	5'd11,	5'd4};
		rom[ 243  ] = { 5'd4,	5'd3,	5'd15,	5'd3};
		rom[ 244  ] = { 5'd8,	5'd0,	5'd8,	5'd19};
		rom[ 245  ] = { 5'd11,	5'd21,	5'd9,	5'd3};
		rom[ 246  ] = { 5'd9,	5'd7,	5'd5,	5'd4};
		rom[ 247  ] = { 5'd10,	5'd7,	5'd5,	5'd4};
		rom[ 248  ] = { 5'd20,	5'd8,	5'd3,	5'd8};
		rom[ 249  ] = { 5'd1,	5'd15,	5'd10,	5'd2};
		rom[ 250  ] = { 5'd14,	5'd17,	5'd10,	5'd2};
		rom[ 251  ] = { 5'd3,	5'd3,	5'd16,	5'd3};
		rom[ 252  ] = { 5'd15,	5'd11,	5'd7,	5'd5};
		rom[ 253  ] = { 5'd11,	5'd1,	5'd2,	5'd13};
		rom[ 254  ] = { 5'd17,	5'd2,	5'd3,	5'd14};
		rom[ 255  ] = { 5'd3,	5'd14,	5'd6,	5'd5};
		rom[ 256  ] = { 5'd7,	5'd8,	5'd10,	5'd2};
		rom[ 257  ] = { 5'd4,	5'd2,	5'd3,	5'd14};
		rom[ 258  ] = { 5'd10,	5'd8,	5'd5,	5'd4};
		rom[ 259  ] = { 5'd8,	5'd17,	5'd8,	5'd5};
		rom[ 260  ] = { 5'd15,	5'd11,	5'd5,	5'd4};
		rom[ 261  ] = { 5'd3,	5'd1,	5'd3,	5'd6};
		rom[ 262  ] = { 5'd12,	5'd16,	5'd6,	5'd3};
		rom[ 263  ] = { 5'd6,	5'd16,	5'd6,	5'd3};
		rom[ 264  ] = { 5'd14,	5'd14,	5'd3,	5'd8};
		rom[ 265  ] = { 5'd1,	5'd14,	5'd13,	5'd2};
		rom[ 266  ] = { 5'd13,	5'd1,	5'd2,	5'd9};
		rom[ 267  ] = { 5'd10,	5'd0,	5'd3,	5'd6};
		rom[ 268  ] = { 5'd12,	5'd2,	5'd3,	5'd9};
		rom[ 269  ] = { 5'd9,	5'd2,	5'd3,	5'd9};
		rom[ 270  ] = { 5'd6,	5'd20,	5'd12,	5'd2};
		rom[ 271  ] = { 5'd9,	5'd6,	5'd2,	5'd9};
		rom[ 272  ] = { 5'd7,	5'd7,	5'd6,	5'd3};
		rom[ 273  ] = { 5'd8,	5'd10,	5'd8,	5'd7};
		rom[ 274  ] = { 5'd7,	5'd8,	5'd10,	5'd4};
		rom[ 275  ] = { 5'd0,	5'd4,	5'd6,	5'd3};
		rom[ 276  ] = { 5'd15,	5'd2,	5'd1,	5'd20};
		rom[ 277  ] = { 5'd0,	5'd6,	5'd6,	5'd3};
		rom[ 278  ] = { 5'd15,	5'd3,	5'd1,	5'd21};
		rom[ 279  ] = { 5'd8,	5'd0,	5'd1,	5'd23};
		rom[ 280  ] = { 5'd15,	5'd10,	5'd9,	5'd2};
		rom[ 281  ] = { 5'd0,	5'd10,	5'd9,	5'd2};
		rom[ 282  ] = { 5'd8,	5'd16,	5'd9,	5'd2};
		rom[ 283  ] = { 5'd0,	5'd16,	5'd9,	5'd2};
		rom[ 284  ] = { 5'd9,	5'd10,	5'd6,	5'd4};
		rom[ 285  ] = { 5'd8,	5'd0,	5'd8,	5'd19};
		rom[ 286  ] = { 5'd9,	5'd7,	5'd8,	5'd6};
		rom[ 287  ] = { 5'd12,	5'd6,	5'd2,	5'd10};
		rom[ 288  ] = { 5'd12,	5'd9,	5'd5,	5'd6};
		rom[ 289  ] = { 5'd6,	5'd0,	5'd1,	5'd19};
		rom[ 290  ] = { 5'd16,	5'd0,	5'd2,	5'd10};
		rom[ 291  ] = { 5'd2,	5'd0,	5'd3,	5'd6};
		rom[ 292  ] = { 5'd0,	5'd12,	5'd24,	5'd1};
		rom[ 293  ] = { 5'd4,	5'd11,	5'd13,	5'd2};
		rom[ 294  ] = { 5'd9,	5'd11,	5'd6,	5'd3};
		rom[ 295  ] = { 5'd0,	5'd14,	5'd16,	5'd2};
		rom[ 296  ] = { 5'd18,	5'd15,	5'd6,	5'd3};
		rom[ 297  ] = { 5'd0,	5'd15,	5'd6,	5'd3};
		rom[ 298  ] = { 5'd8,	5'd7,	5'd5,	5'd4};
		rom[ 299  ] = { 5'd10,	5'd7,	5'd2,	5'd9};
		rom[ 300  ] = { 5'd13,	5'd0,	5'd2,	5'd9};
		rom[ 301  ] = { 5'd9,	5'd0,	5'd2,	5'd9};
		rom[ 302  ] = { 5'd14,	5'd3,	5'd2,	5'd15};
		rom[ 303  ] = { 5'd8,	5'd3,	5'd2,	5'd15};
		rom[ 304  ] = { 5'd15,	5'd4,	5'd9,	5'd2};
		rom[ 305  ] = { 5'd8,	5'd10,	5'd3,	5'd7};
		rom[ 306  ] = { 5'd9,	5'd19,	5'd6,	5'd5};
		rom[ 307  ] = { 5'd7,	5'd17,	5'd5,	5'd4};
		rom[ 308  ] = { 5'd14,	5'd13,	5'd3,	5'd8};
		rom[ 309  ] = { 5'd2,	5'd18,	5'd18,	5'd1};
		rom[ 310  ] = { 5'd5,	5'd19,	5'd19,	5'd1};
		rom[ 311  ] = { 5'd11,	5'd0,	5'd2,	5'd9};
		rom[ 312  ] = { 5'd13,	5'd4,	5'd1,	5'd18};
		rom[ 313  ] = { 5'd10,	5'd4,	5'd1,	5'd18};
		rom[ 314  ] = { 5'd9,	5'd3,	5'd6,	5'd9};
		rom[ 315  ] = { 5'd8,	5'd1,	5'd2,	5'd14};
		rom[ 316  ] = { 5'd12,	5'd19,	5'd9,	5'd3};
		rom[ 317  ] = { 5'd1,	5'd3,	5'd10,	5'd8};
		rom[ 318  ] = { 5'd15,	5'd5,	5'd3,	5'd6};
		rom[ 319  ] = { 5'd1,	5'd2,	5'd11,	5'd8};
		rom[ 320  ] = { 5'd10,	5'd19,	5'd5,	5'd5};
		rom[ 321  ] = { 5'd3,	5'd22,	5'd18,	5'd1};
		rom[ 322  ] = { 5'd12,	5'd14,	5'd2,	5'd10};
		rom[ 323  ] = { 5'd8,	5'd2,	5'd8,	5'd4};
		rom[ 324  ] = { 5'd6,	5'd7,	5'd12,	5'd3};
		rom[ 325  ] = { 5'd10,	5'd6,	5'd4,	5'd5};
		rom[ 326  ] = { 5'd5,	5'd12,	5'd14,	5'd4};
		rom[ 327  ] = { 5'd4,	5'd14,	5'd4,	5'd5};
		rom[ 328  ] = { 5'd11,	5'd13,	5'd5,	5'd7};
		rom[ 329  ] = { 5'd7,	5'd14,	5'd3,	5'd8};
		rom[ 330  ] = { 5'd9,	5'd7,	5'd6,	5'd8};
		rom[ 331  ] = { 5'd2,	5'd4,	5'd20,	5'd1};
		rom[ 332  ] = { 5'd3,	5'd14,	5'd19,	5'd2};
		rom[ 333  ] = { 5'd10,	5'd6,	5'd2,	5'd9};
		rom[ 334  ] = { 5'd16,	5'd6,	5'd3,	5'd14};
		rom[ 335  ] = { 5'd9,	5'd9,	5'd2,	5'd12};
		rom[ 336  ] = { 5'd21,	5'd6,	5'd3,	5'd9};
		rom[ 337  ] = { 5'd0,	5'd6,	5'd3,	5'd9};
		rom[ 338  ] = { 5'd18,	5'd5,	5'd6,	5'd3};
		rom[ 339  ] = { 5'd3,	5'd20,	5'd15,	5'd2};
		rom[ 340  ] = { 5'd18,	5'd5,	5'd6,	5'd3};
		rom[ 341  ] = { 5'd0,	5'd5,	5'd6,	5'd3};
		rom[ 342  ] = { 5'd5,	5'd11,	5'd18,	5'd1};
		rom[ 343  ] = { 5'd6,	5'd2,	5'd12,	5'd2};
		rom[ 344  ] = { 5'd12,	5'd0,	5'd2,	5'd9};
		rom[ 345  ] = { 5'd10,	5'd0,	5'd2,	5'd9};
		rom[ 346  ] = { 5'd15,	5'd14,	5'd9,	5'd2};
		rom[ 347  ] = { 5'd3,	5'd8,	5'd13,	5'd2};
		rom[ 348  ] = { 5'd15,	5'd14,	5'd9,	5'd2};
		rom[ 349  ] = { 5'd5,	5'd5,	5'd3,	5'd15};
		rom[ 350  ] = { 5'd11,	5'd8,	5'd3,	5'd6};
		rom[ 351  ] = { 5'd8,	5'd13,	5'd3,	5'd7};
		rom[ 352  ] = { 5'd15,	5'd14,	5'd9,	5'd2};
		rom[ 353  ] = { 5'd9,	5'd12,	5'd5,	5'd4};
		rom[ 354  ] = { 5'd13,	5'd1,	5'd2,	5'd19};
		rom[ 355  ] = { 5'd9,	5'd1,	5'd2,	5'd19};
		rom[ 356  ] = { 5'd18,	5'd12,	5'd6,	5'd3};
		rom[ 357  ] = { 5'd1,	5'd22,	5'd18,	5'd1};
		rom[ 358  ] = { 5'd14,	5'd16,	5'd10,	5'd3};
		rom[ 359  ] = { 5'd1,	5'd13,	5'd11,	5'd2};
		rom[ 360  ] = { 5'd12,	5'd6,	5'd8,	5'd3};
		rom[ 361  ] = { 5'd1,	5'd0,	5'd9,	5'd11};
		rom[ 362  ] = { 5'd14,	5'd7,	5'd4,	5'd7};
		rom[ 363  ] = { 5'd0,	5'd4,	5'd3,	5'd10};
		rom[ 364  ] = { 5'd17,	5'd0,	5'd2,	5'd9};
		rom[ 365  ] = { 5'd5,	5'd0,	5'd2,	5'd9};
		rom[ 366  ] = { 5'd18,	5'd12,	5'd3,	5'd6};
		rom[ 367  ] = { 5'd3,	5'd12,	5'd3,	5'd6};
		rom[ 368  ] = { 5'd15,	5'd14,	5'd9,	5'd2};
		rom[ 369  ] = { 5'd0,	5'd14,	5'd9,	5'd2};
		rom[ 370  ] = { 5'd4,	5'd15,	5'd19,	5'd1};
		rom[ 371  ] = { 5'd2,	5'd14,	5'd19,	5'd1};
		rom[ 372  ] = { 5'd14,	5'd17,	5'd10,	5'd2};
		rom[ 373  ] = { 5'd6,	5'd0,	5'd5,	5'd6};
		rom[ 374  ] = { 5'd20,	5'd1,	5'd3,	5'd6};
		rom[ 375  ] = { 5'd1,	5'd1,	5'd3,	5'd6};
		rom[ 376  ] = { 5'd16,	5'd17,	5'd6,	5'd3};
		rom[ 377  ] = { 5'd7,	5'd9,	5'd9,	5'd6};
		rom[ 378  ] = { 5'd12,	5'd7,	5'd4,	5'd6};
		rom[ 379  ] = { 5'd4,	5'd4,	5'd14,	5'd4};
		rom[ 380  ] = { 5'd12,	5'd6,	5'd2,	5'd9};
		rom[ 381  ] = { 5'd8,	5'd10,	5'd6,	5'd3};
		rom[ 382  ] = { 5'd15,	5'd17,	5'd9,	5'd2};
		rom[ 383  ] = { 5'd7,	5'd1,	5'd7,	5'd23};
		rom[ 384  ] = { 5'd6,	5'd11,	5'd17,	5'd2};
		rom[ 385  ] = { 5'd1,	5'd6,	5'd11,	5'd6};
		rom[ 386  ] = { 5'd6,	5'd17,	5'd13,	5'd2};
		rom[ 387  ] = { 5'd0,	5'd17,	5'd9,	5'd2};
		rom[ 388  ] = { 5'd13,	5'd7,	5'd5,	5'd4};
		rom[ 389  ] = { 5'd9,	5'd15,	5'd6,	5'd3};
		rom[ 390  ] = { 5'd12,	5'd8,	5'd6,	5'd3};
		rom[ 391  ] = { 5'd8,	5'd14,	5'd8,	5'd4};
		rom[ 392  ] = { 5'd16,	5'd16,	5'd3,	5'd6};
		rom[ 393  ] = { 5'd0,	5'd4,	5'd24,	5'd1};
		rom[ 394  ] = { 5'd14,	5'd19,	5'd10,	5'd2};
		rom[ 395  ] = { 5'd7,	5'd13,	5'd6,	5'd3};
		rom[ 396  ] = { 5'd5,	5'd3,	5'd18,	5'd3};
		rom[ 397  ] = { 5'd4,	5'd6,	5'd16,	5'd3};
		rom[ 398  ] = { 5'd16,	5'd11,	5'd3,	5'd6};
		rom[ 399  ] = { 5'd6,	5'd7,	5'd6,	5'd4};
		rom[ 400  ] = { 5'd12,	5'd6,	5'd2,	5'd9};
		rom[ 401  ] = { 5'd11,	5'd8,	5'd2,	5'd10};
		rom[ 402  ] = { 5'd11,	5'd15,	5'd2,	5'd9};
		rom[ 403  ] = { 5'd12,	5'd1,	5'd9,	5'd21};
		rom[ 404  ] = { 5'd6,	5'd8,	5'd6,	5'd7};
		rom[ 405  ] = { 5'd10,	5'd5,	5'd2,	5'd9};
		rom[ 406  ] = { 5'd8,	5'd2,	5'd8,	5'd4};
		rom[ 407  ] = { 5'd14,	5'd11,	5'd5,	5'd4};
		rom[ 408  ] = { 5'd5,	5'd11,	5'd5,	5'd4};
		rom[ 409  ] = { 5'd11,	5'd6,	5'd2,	5'd9};
		rom[ 410  ] = { 5'd3,	5'd1,	5'd3,	5'd17};
		rom[ 411  ] = { 5'd3,	5'd4,	5'd19,	5'd3};
		rom[ 412  ] = { 5'd3,	5'd18,	5'd6,	5'd3};
		rom[ 413  ] = { 5'd20,	5'd4,	5'd2,	5'd19};
		rom[ 414  ] = { 5'd5,	5'd16,	5'd5,	5'd7};
		rom[ 415  ] = { 5'd13,	5'd7,	5'd5,	5'd6};
		rom[ 416  ] = { 5'd6,	5'd7,	5'd5,	5'd6};
		rom[ 417  ] = { 5'd12,	5'd2,	5'd3,	5'd6};
		rom[ 418  ] = { 5'd8,	5'd20,	5'd7,	5'd4};
		rom[ 419  ] = { 5'd9,	5'd14,	5'd9,	5'd2};
		rom[ 420  ] = { 5'd10,	5'd2,	5'd3,	5'd6};
		rom[ 421  ] = { 5'd13,	5'd0,	5'd2,	5'd14};
		rom[ 422  ] = { 5'd9,	5'd0,	5'd2,	5'd14};
		rom[ 423  ] = { 5'd14,	5'd17,	5'd9,	5'd2};
		rom[ 424  ] = { 5'd8,	5'd8,	5'd6,	5'd5};
		rom[ 425  ] = { 5'd20,	5'd3,	5'd2,	5'd11};
		rom[ 426  ] = { 5'd6,	5'd12,	5'd11,	5'd7};
		rom[ 427  ] = { 5'd18,	5'd7,	5'd6,	5'd3};
		rom[ 428  ] = { 5'd7,	5'd8,	5'd9,	5'd2};
		rom[ 429  ] = { 5'd18,	5'd7,	5'd6,	5'd3};
		rom[ 430  ] = { 5'd0,	5'd7,	5'd6,	5'd3};
		rom[ 431  ] = { 5'd9,	5'd6,	5'd9,	5'd2};
		rom[ 432  ] = { 5'd0,	5'd23,	5'd19,	5'd1};
		rom[ 433  ] = { 5'd17,	5'd17,	5'd6,	5'd3};
		rom[ 434  ] = { 5'd1,	5'd17,	5'd6,	5'd3};
		rom[ 435  ] = { 5'd14,	5'd11,	5'd2,	5'd9};
		rom[ 436  ] = { 5'd8,	5'd11,	5'd2,	5'd9};
		rom[ 437  ] = { 5'd9,	5'd9,	5'd6,	5'd7};
		rom[ 438  ] = { 5'd9,	5'd17,	5'd6,	5'd5};
		rom[ 439  ] = { 5'd14,	5'd0,	5'd2,	5'd9};
		rom[ 440  ] = { 5'd8,	5'd0,	5'd2,	5'd9};
		rom[ 441  ] = { 5'd6,	5'd18,	5'd18,	5'd1};
		rom[ 442  ] = { 5'd1,	5'd18,	5'd18,	5'd1};
		rom[ 443  ] = { 5'd10,	5'd12,	5'd11,	5'd6};
		rom[ 444  ] = { 5'd5,	5'd6,	5'd7,	5'd3};
		rom[ 445  ] = { 5'd5,	5'd6,	5'd15,	5'd2};
		rom[ 446  ] = { 5'd0,	5'd1,	5'd22,	5'd1};
		rom[ 447  ] = { 5'd8,	5'd0,	5'd8,	5'd24};
		rom[ 448  ] = { 5'd10,	5'd15,	5'd9,	5'd4};
		rom[ 449  ] = { 5'd6,	5'd11,	5'd12,	5'd3};
		rom[ 450  ] = { 5'd4,	5'd16,	5'd7,	5'd4};
		rom[ 451  ] = { 5'd12,	5'd2,	5'd11,	5'd3};
		rom[ 452  ] = { 5'd12,	5'd20,	5'd7,	5'd3};
		rom[ 453  ] = { 5'd12,	5'd0,	5'd12,	5'd8};
		rom[ 454  ] = { 5'd3,	5'd13,	5'd9,	5'd2};
		rom[ 455  ] = { 5'd2,	5'd11,	5'd22,	5'd1};
		rom[ 456  ] = { 5'd6,	5'd7,	5'd11,	5'd4};
		rom[ 457  ] = { 5'd14,	5'd8,	5'd6,	5'd3};
		rom[ 458  ] = { 5'd0,	5'd9,	5'd24,	5'd2};
		rom[ 459  ] = { 5'd19,	5'd0,	5'd5,	5'd5};
		rom[ 460  ] = { 5'd0,	5'd0,	5'd5,	5'd5};
		rom[ 461  ] = { 5'd12,	5'd1,	5'd12,	5'd2};
		rom[ 462  ] = { 5'd0,	5'd18,	5'd18,	5'd1};
		rom[ 463  ] = { 5'd13,	5'd15,	5'd8,	5'd3};
		rom[ 464  ] = { 5'd3,	5'd15,	5'd8,	5'd3};
		rom[ 465  ] = { 5'd6,	5'd17,	5'd18,	5'd1};
		rom[ 466  ] = { 5'd0,	5'd18,	5'd21,	5'd5};
		rom[ 467  ] = { 5'd15,	5'd0,	5'd2,	5'd24};
		rom[ 468  ] = { 5'd9,	5'd4,	5'd2,	5'd11};
		rom[ 469  ] = { 5'd12,	5'd5,	5'd3,	5'd6};
		rom[ 470  ] = { 5'd1,	5'd14,	5'd2,	5'd10};
		rom[ 471  ] = { 5'd15,	5'd0,	5'd2,	5'd24};
		rom[ 472  ] = { 5'd7,	5'd0,	5'd2,	5'd24};
		rom[ 473  ] = { 5'd19,	5'd7,	5'd3,	5'd7};
		rom[ 474  ] = { 5'd6,	5'd7,	5'd2,	5'd12};
		rom[ 475  ] = { 5'd8,	5'd5,	5'd8,	5'd14};
		rom[ 476  ] = { 5'd5,	5'd15,	5'd10,	5'd2};
		rom[ 477  ] = { 5'd14,	5'd0,	5'd2,	5'd9};
		rom[ 478  ] = { 5'd2,	5'd7,	5'd3,	5'd7};
		rom[ 479  ] = { 5'd18,	5'd2,	5'd3,	5'd15};
		rom[ 480  ] = { 5'd2,	5'd2,	5'd2,	5'd9};
		rom[ 481  ] = { 5'd17,	5'd2,	5'd5,	5'd7};
		rom[ 482  ] = { 5'd12,	5'd6,	5'd1,	5'd18};
		rom[ 483  ] = { 5'd14,	5'd5,	5'd5,	5'd6};
		rom[ 484  ] = { 5'd10,	5'd6,	5'd2,	5'd10};
		rom[ 485  ] = { 5'd14,	5'd0,	5'd2,	5'd9};
		rom[ 486  ] = { 5'd6,	5'd3,	5'd3,	5'd7};
		rom[ 487  ] = { 5'd6,	5'd7,	5'd7,	5'd3};
		rom[ 488  ] = { 5'd11,	5'd7,	5'd4,	5'd6};
		rom[ 489  ] = { 5'd12,	5'd13,	5'd7,	5'd6};
		rom[ 490  ] = { 5'd10,	5'd6,	5'd2,	5'd9};
		rom[ 491  ] = { 5'd16,	5'd17,	5'd6,	5'd3};
		rom[ 492  ] = { 5'd6,	5'd0,	5'd2,	5'd13};
		rom[ 493  ] = { 5'd9,	5'd2,	5'd7,	5'd3};
		rom[ 494  ] = { 5'd5,	5'd8,	5'd5,	5'd4};
		rom[ 495  ] = { 5'd10,	5'd8,	5'd4,	5'd5};
		rom[ 496  ] = { 5'd8,	5'd8,	5'd5,	5'd4};
		rom[ 497  ] = { 5'd6,	5'd3,	5'd11,	5'd3};
		rom[ 498  ] = { 5'd10,	5'd6,	5'd4,	5'd5};
		rom[ 499  ] = { 5'd8,	5'd0,	5'd8,	5'd5};
		rom[ 500  ] = { 5'd1,	5'd12,	5'd23,	5'd2};
		rom[ 501  ] = { 5'd9,	5'd21,	5'd6,	5'd3};
		rom[ 502  ] = { 5'd3,	5'd8,	5'd21,	5'd2};
		rom[ 503  ] = { 5'd2,	5'd5,	5'd2,	5'd12};
		rom[ 504  ] = { 5'd10,	5'd7,	5'd4,	5'd5};
		rom[ 505  ] = { 5'd8,	5'd12,	5'd8,	5'd5};
		rom[ 506  ] = { 5'd10,	5'd7,	5'd5,	5'd12};
		rom[ 507  ] = { 5'd0,	5'd19,	5'd10,	5'd2};
		rom[ 508  ] = { 5'd14,	5'd20,	5'd9,	5'd2};
		rom[ 509  ] = { 5'd9,	5'd14,	5'd6,	5'd8};
		rom[ 510  ] = { 5'd14,	5'd20,	5'd9,	5'd2};
		rom[ 511  ] = { 5'd1,	5'd20,	5'd9,	5'd2};
		rom[ 512  ] = { 5'd15,	5'd11,	5'd9,	5'd2};
		rom[ 513  ] = { 5'd0,	5'd11,	5'd9,	5'd2};
		rom[ 514  ] = { 5'd19,	5'd3,	5'd2,	5'd9};
		rom[ 515  ] = { 5'd2,	5'd18,	5'd18,	5'd1};
		rom[ 516  ] = { 5'd3,	5'd17,	5'd21,	5'd2};
		rom[ 517  ] = { 5'd9,	5'd20,	5'd6,	5'd3};
		rom[ 518  ] = { 5'd18,	5'd6,	5'd6,	5'd3};
		rom[ 519  ] = { 5'd0,	5'd6,	5'd6,	5'd3};
		rom[ 520  ] = { 5'd12,	5'd0,	5'd8,	5'd5};
		rom[ 521  ] = { 5'd2,	5'd0,	5'd5,	5'd8};
		rom[ 522  ] = { 5'd14,	5'd0,	5'd5,	5'd5};
		rom[ 523  ] = { 5'd5,	5'd0,	5'd5,	5'd5};
		rom[ 524  ] = { 5'd18,	5'd3,	5'd3,	5'd10};
		rom[ 525  ] = { 5'd5,	5'd11,	5'd6,	5'd3};
		rom[ 526  ] = { 5'd22,	5'd0,	5'd1,	5'd18};
		rom[ 527  ] = { 5'd8,	5'd0,	5'd2,	5'd9};
		rom[ 528  ] = { 5'd11,	5'd8,	5'd3,	5'd7};
		rom[ 529  ] = { 5'd7,	5'd12,	5'd4,	5'd5};
		rom[ 530  ] = { 5'd22,	5'd0,	5'd1,	5'd18};
		rom[ 531  ] = { 5'd12,	5'd6,	5'd2,	5'd9};
		rom[ 532  ] = { 5'd15,	5'd2,	5'd9,	5'd2};
		rom[ 533  ] = { 5'd0,	5'd3,	5'd24,	5'd1};
		rom[ 534  ] = { 5'd13,	5'd7,	5'd2,	5'd9};
		rom[ 535  ] = { 5'd9,	5'd6,	5'd2,	5'd10};
		rom[ 536  ] = { 5'd14,	5'd1,	5'd2,	5'd12};
		rom[ 537  ] = { 5'd6,	5'd10,	5'd12,	5'd6};
		rom[ 538  ] = { 5'd14,	5'd3,	5'd1,	5'd21};
		rom[ 539  ] = { 5'd6,	5'd5,	5'd12,	5'd4};
		rom[ 540  ] = { 5'd3,	5'd4,	5'd18,	5'd4};
		rom[ 541  ] = { 5'd3,	5'd1,	5'd18,	5'd1};
		rom[ 542  ] = { 5'd12,	5'd13,	5'd12,	5'd2};
		rom[ 543  ] = { 5'd12,	5'd5,	5'd2,	5'd9};
		rom[ 544  ] = { 5'd13,	5'd1,	5'd2,	5'd9};
		rom[ 545  ] = { 5'd8,	5'd2,	5'd2,	5'd22};
		rom[ 546  ] = { 5'd20,	5'd10,	5'd4,	5'd7};
		rom[ 547  ] = { 5'd3,	5'd9,	5'd16,	5'd5};
		rom[ 548  ] = { 5'd20,	5'd10,	5'd4,	5'd7};
		rom[ 549  ] = { 5'd0,	5'd10,	5'd4,	5'd7};
		rom[ 550  ] = { 5'd10,	5'd17,	5'd11,	5'd3};
		rom[ 551  ] = { 5'd8,	5'd7,	5'd8,	5'd9};
		rom[ 552  ] = { 5'd13,	5'd1,	5'd2,	5'd16};
		rom[ 553  ] = { 5'd9,	5'd1,	5'd2,	5'd16};
		rom[ 554  ] = { 5'd13,	5'd5,	5'd8,	5'd4};
		rom[ 555  ] = { 5'd0,	5'd12,	5'd6,	5'd3};
		rom[ 556  ] = { 5'd6,	5'd17,	5'd18,	5'd1};
		rom[ 557  ] = { 5'd3,	5'd15,	5'd6,	5'd3};
		rom[ 558  ] = { 5'd8,	5'd16,	5'd9,	5'd2};
		rom[ 559  ] = { 5'd2,	5'd13,	5'd4,	5'd5};
		rom[ 560  ] = { 5'd15,	5'd11,	5'd3,	5'd6};
		rom[ 561  ] = { 5'd3,	5'd6,	5'd18,	5'd1};
		rom[ 562  ] = { 5'd19,	5'd5,	5'd2,	5'd11};
		rom[ 563  ] = { 5'd3,	5'd5,	5'd2,	5'd11};
		rom[ 564  ] = { 5'd19,	5'd1,	5'd2,	5'd9};
		rom[ 565  ] = { 5'd3,	5'd1,	5'd2,	5'd9};
		rom[ 566  ] = { 5'd4,	5'd15,	5'd9,	5'd9};
		rom[ 567  ] = { 5'd6,	5'd11,	5'd12,	5'd2};
		rom[ 568  ] = { 5'd15,	5'd4,	5'd9,	5'd2};
		rom[ 569  ] = { 5'd0,	5'd4,	5'd9,	5'd2};
		rom[ 570  ] = { 5'd17,	5'd0,	5'd2,	5'd17};
		rom[ 571  ] = { 5'd5,	5'd0,	5'd2,	5'd17};
		rom[ 572  ] = { 5'd8,	5'd19,	5'd9,	5'd2};
		rom[ 573  ] = { 5'd6,	5'd11,	5'd3,	5'd6};
		rom[ 574  ] = { 5'd5,	5'd8,	5'd14,	5'd6};
		rom[ 575  ] = { 5'd10,	5'd8,	5'd3,	5'd6};
		rom[ 576  ] = { 5'd10,	5'd12,	5'd14,	5'd5};
		rom[ 577  ] = { 5'd0,	5'd12,	5'd14,	5'd5};
		rom[ 578  ] = { 5'd15,	5'd2,	5'd9,	5'd2};
		rom[ 579  ] = { 5'd0,	5'd2,	5'd9,	5'd2};
		rom[ 580  ] = { 5'd14,	5'd6,	5'd2,	5'd14};
		rom[ 581  ] = { 5'd11,	5'd7,	5'd2,	5'd9};
		rom[ 582  ] = { 5'd14,	5'd6,	5'd2,	5'd15};
		rom[ 583  ] = { 5'd8,	5'd6,	5'd2,	5'd15};
		rom[ 584  ] = { 5'd15,	5'd3,	5'd4,	5'd9};
		rom[ 585  ] = { 5'd3,	5'd0,	5'd3,	5'd21};
		rom[ 586  ] = { 5'd11,	5'd13,	5'd8,	5'd4};
		rom[ 587  ] = { 5'd6,	5'd7,	5'd5,	5'd6};
		rom[ 588  ] = { 5'd12,	5'd6,	5'd2,	5'd9};
		rom[ 589  ] = { 5'd0,	5'd3,	5'd6,	5'd3};
		rom[ 590  ] = { 5'd3,	5'd15,	5'd18,	5'd1};
		rom[ 591  ] = { 5'd3,	5'd14,	5'd4,	5'd5};
		rom[ 592  ] = { 5'd12,	5'd12,	5'd12,	5'd2};
		rom[ 593  ] = { 5'd1,	5'd2,	5'd1,	5'd20};
		rom[ 594  ] = { 5'd17,	5'd16,	5'd5,	5'd4};
		rom[ 595  ] = { 5'd2,	5'd16,	5'd5,	5'd4};
		rom[ 596  ] = { 5'd7,	5'd3,	5'd10,	5'd3};
		rom[ 597  ] = { 5'd8,	5'd0,	5'd8,	5'd3};
		rom[ 598  ] = { 5'd3,	5'd10,	5'd15,	5'd2};
		rom[ 599  ] = { 5'd10,	5'd5,	5'd4,	5'd6};
		rom[ 600  ] = { 5'd5,	5'd16,	5'd14,	5'd3};
		rom[ 601  ] = { 5'd11,	5'd19,	5'd4,	5'd5};
		rom[ 602  ] = { 5'd3,	5'd6,	5'd3,	5'd7};
		rom[ 603  ] = { 5'd18,	5'd0,	5'd3,	5'd6};
		rom[ 604  ] = { 5'd3,	5'd2,	5'd18,	5'd1};
		rom[ 605  ] = { 5'd9,	5'd12,	5'd14,	5'd6};
		rom[ 606  ] = { 5'd3,	5'd0,	5'd3,	5'd6};
		rom[ 607  ] = { 5'd13,	5'd11,	5'd3,	5'd6};
		rom[ 608  ] = { 5'd8,	5'd20,	5'd8,	5'd3};
		rom[ 609  ] = { 5'd13,	5'd11,	5'd3,	5'd7};
		rom[ 610  ] = { 5'd4,	5'd14,	5'd10,	5'd2};
		rom[ 611  ] = { 5'd13,	5'd11,	5'd3,	5'd6};
		rom[ 612  ] = { 5'd8,	5'd11,	5'd3,	5'd7};
		rom[ 613  ] = { 5'd7,	5'd8,	5'd11,	5'd4};
		rom[ 614  ] = { 5'd6,	5'd17,	5'd10,	5'd2};
		rom[ 615  ] = { 5'd16,	5'd0,	5'd2,	5'd9};
		rom[ 616  ] = { 5'd6,	5'd0,	5'd2,	5'd9};
		rom[ 617  ] = { 5'd11,	5'd7,	5'd4,	5'd5};
		rom[ 618  ] = { 5'd0,	5'd1,	5'd20,	5'd1};
		rom[ 619  ] = { 5'd13,	5'd20,	5'd10,	5'd2};
		rom[ 620  ] = { 5'd5,	5'd7,	5'd3,	5'd11};
		rom[ 621  ] = { 5'd10,	5'd17,	5'd10,	5'd3};
		rom[ 622  ] = { 5'd10,	5'd2,	5'd2,	5'd9};
		rom[ 623  ] = { 5'd14,	5'd3,	5'd5,	5'd4};
		rom[ 624  ] = { 5'd6,	5'd6,	5'd6,	5'd3};
		rom[ 625  ] = { 5'd12,	5'd8,	5'd4,	5'd5};
		rom[ 626  ] = { 5'd7,	5'd12,	5'd4,	5'd8};
		rom[ 627  ] = { 5'd8,	5'd10,	5'd9,	5'd2};
		rom[ 628  ] = { 5'd5,	5'd5,	5'd14,	5'd3};
		rom[ 629  ] = { 5'd3,	5'd20,	5'd19,	5'd4};
		rom[ 630  ] = { 5'd5,	5'd0,	5'd5,	5'd8};
		rom[ 631  ] = { 5'd5,	5'd2,	5'd8,	5'd18};
		rom[ 632  ] = { 5'd8,	5'd11,	5'd8,	5'd11};
		rom[ 633  ] = { 5'd3,	5'd3,	5'd9,	5'd5};
		rom[ 634  ] = { 5'd1,	5'd17,	5'd18,	5'd1};
		rom[ 635  ] = { 5'd5,	5'd18,	5'd18,	5'd1};
		rom[ 636  ] = { 5'd1,	5'd15,	5'd9,	5'd2};
		rom[ 637  ] = { 5'd1,	5'd14,	5'd23,	5'd5};
		rom[ 638  ] = { 5'd3,	5'd8,	5'd18,	5'd1};
		rom[ 639  ] = { 5'd6,	5'd8,	5'd6,	5'd3};
		rom[ 640  ] = { 5'd7,	5'd2,	5'd1,	5'd22};
		rom[ 641  ] = { 5'd14,	5'd19,	5'd10,	5'd2};
		rom[ 642  ] = { 5'd1,	5'd20,	5'd10,	5'd2};
		rom[ 643  ] = { 5'd13,	5'd3,	5'd2,	5'd12};
		rom[ 644  ] = { 5'd12,	5'd6,	5'd2,	5'd9};
		rom[ 645  ] = { 5'd13,	5'd0,	5'd2,	5'd9};
		rom[ 646  ] = { 5'd9,	5'd0,	5'd2,	5'd9};
		rom[ 647  ] = { 5'd15,	5'd10,	5'd3,	5'd6};
		rom[ 648  ] = { 5'd5,	5'd11,	5'd3,	5'd9};
		rom[ 649  ] = { 5'd15,	5'd5,	5'd1,	5'd19};
		rom[ 650  ] = { 5'd6,	5'd8,	5'd9,	5'd2};
		rom[ 651  ] = { 5'd15,	5'd5,	5'd1,	5'd19};
		rom[ 652  ] = { 5'd0,	5'd6,	5'd6,	5'd3};
		rom[ 653  ] = { 5'd5,	5'd22,	5'd18,	5'd1};
		rom[ 654  ] = { 5'd7,	5'd10,	5'd6,	5'd4};
		rom[ 655  ] = { 5'd17,	5'd4,	5'd4,	5'd5};
		rom[ 656  ] = { 5'd10,	5'd8,	5'd3,	5'd6};
		rom[ 657  ] = { 5'd15,	5'd9,	5'd3,	5'd8};
		rom[ 658  ] = { 5'd0,	5'd10,	5'd5,	5'd4};
		rom[ 659  ] = { 5'd14,	5'd6,	5'd7,	5'd3};
		rom[ 660  ] = { 5'd8,	5'd5,	5'd1,	5'd19};
		rom[ 661  ] = { 5'd13,	5'd4,	5'd5,	5'd20};
		rom[ 662  ] = { 5'd6,	5'd4,	5'd5,	5'd20};
		rom[ 663  ] = { 5'd13,	5'd10,	5'd3,	5'd6};
		rom[ 664  ] = { 5'd8,	5'd10,	5'd3,	5'd6};
		rom[ 665  ] = { 5'd17,	5'd2,	5'd3,	5'd7};
		rom[ 666  ] = { 5'd4,	5'd2,	5'd3,	5'd7};
		rom[ 667  ] = { 5'd12,	5'd4,	5'd3,	5'd7};
		rom[ 668  ] = { 5'd11,	5'd4,	5'd2,	5'd9};
		rom[ 669  ] = { 5'd11,	5'd4,	5'd4,	5'd10};
		rom[ 670  ] = { 5'd9,	5'd4,	5'd4,	5'd10};
		rom[ 671  ] = { 5'd8,	5'd20,	5'd10,	5'd2};
		rom[ 672  ] = { 5'd1,	5'd20,	5'd21,	5'd2};
		rom[ 673  ] = { 5'd9,	5'd2,	5'd6,	5'd6};
		rom[ 674  ] = { 5'd9,	5'd2,	5'd6,	5'd6};
		rom[ 675  ] = { 5'd18,	5'd5,	5'd6,	5'd3};
		rom[ 676  ] = { 5'd8,	5'd11,	5'd6,	5'd3};
		rom[ 677  ] = { 5'd2,	5'd9,	5'd20,	5'd2};
		rom[ 678  ] = { 5'd0,	5'd5,	5'd6,	5'd3};
		rom[ 679  ] = { 5'd18,	5'd14,	5'd4,	5'd5};
		rom[ 680  ] = { 5'd2,	5'd14,	5'd4,	5'd5};
		rom[ 681  ] = { 5'd2,	5'd11,	5'd10,	5'd13};
		rom[ 682  ] = { 5'd12,	5'd9,	5'd6,	5'd5};
		rom[ 683  ] = { 5'd13,	5'd6,	5'd8,	5'd3};
		rom[ 684  ] = { 5'd1,	5'd21,	5'd9,	5'd2};
		rom[ 685  ] = { 5'd11,	5'd5,	5'd4,	5'd5};
		rom[ 686  ] = { 5'd3,	5'd5,	5'd7,	5'd6};
		rom[ 687  ] = { 5'd12,	5'd4,	5'd3,	5'd6};
		rom[ 688  ] = { 5'd2,	5'd7,	5'd19,	5'd1};
		rom[ 689  ] = { 5'd18,	5'd13,	5'd6,	5'd3};
		rom[ 690  ] = { 5'd3,	5'd8,	5'd18,	5'd1};
		rom[ 691  ] = { 5'd22,	5'd2,	5'd2,	5'd9};
		rom[ 692  ] = { 5'd2,	5'd19,	5'd20,	5'd1};
		rom[ 693  ] = { 5'd1,	5'd10,	5'd22,	5'd1};
		rom[ 694  ] = { 5'd0,	5'd2,	5'd2,	5'd9};
		rom[ 695  ] = { 5'd19,	5'd0,	5'd2,	5'd23};
		rom[ 696  ] = { 5'd3,	5'd3,	5'd3,	5'd19};
		rom[ 697  ] = { 5'd20,	5'd2,	5'd2,	5'd9};
		rom[ 698  ] = { 5'd0,	5'd7,	5'd10,	5'd2};
		rom[ 699  ] = { 5'd13,	5'd0,	5'd6,	5'd6};
		rom[ 700  ] = { 5'd0,	5'd3,	5'd12,	5'd3};
		rom[ 701  ] = { 5'd10,	5'd19,	5'd4,	5'd5};
		rom[ 702  ] = { 5'd8,	5'd14,	5'd4,	5'd5};
		rom[ 703  ] = { 5'd4,	5'd14,	5'd17,	5'd3};
		rom[ 704  ] = { 5'd2,	5'd5,	5'd9,	5'd4};
		rom[ 705  ] = { 5'd14,	5'd6,	5'd7,	5'd3};
		rom[ 706  ] = { 5'd3,	5'd6,	5'd7,	5'd3};
		rom[ 707  ] = { 5'd17,	5'd5,	5'd1,	5'd18};
		rom[ 708  ] = { 5'd6,	5'd5,	5'd1,	5'd18};
		rom[ 709  ] = { 5'd10,	5'd12,	5'd14,	5'd2};
		rom[ 710  ] = { 5'd4,	5'd12,	5'd9,	5'd2};
		rom[ 711  ] = { 5'd2,	5'd3,	5'd18,	5'd3};
		rom[ 712  ] = { 5'd10,	5'd3,	5'd4,	5'd8};
		rom[ 713  ] = { 5'd5,	5'd1,	5'd4,	5'd5};
		rom[ 714  ] = { 5'd12,	5'd11,	5'd7,	5'd4};
		rom[ 715  ] = { 5'd0,	5'd14,	5'd22,	5'd2};
		rom[ 716  ] = { 5'd15,	5'd11,	5'd4,	5'd5};
		rom[ 717  ] = { 5'd5,	5'd11,	5'd7,	5'd4};
		rom[ 718  ] = { 5'd8,	5'd20,	5'd9,	5'd2};
		rom[ 719  ] = { 5'd1,	5'd4,	5'd22,	5'd2};
		rom[ 720  ] = { 5'd19,	5'd3,	5'd2,	5'd17};
		rom[ 721  ] = { 5'd8,	5'd11,	5'd8,	5'd9};
		rom[ 722  ] = { 5'd20,	5'd0,	5'd3,	5'd6};
		rom[ 723  ] = { 5'd9,	5'd0,	5'd2,	5'd9};
		rom[ 724  ] = { 5'd15,	5'd11,	5'd9,	5'd6};
		rom[ 725  ] = { 5'd2,	5'd23,	5'd18,	5'd1};
		rom[ 726  ] = { 5'd16,	5'd10,	5'd6,	5'd3};
		rom[ 727  ] = { 5'd2,	5'd1,	5'd2,	5'd11};
		rom[ 728  ] = { 5'd20,	5'd0,	5'd2,	5'd10};
		rom[ 729  ] = { 5'd3,	5'd3,	5'd2,	5'd17};
		rom[ 730  ] = { 5'd15,	5'd17,	5'd9,	5'd2};
		rom[ 731  ] = { 5'd0,	5'd16,	5'd8,	5'd3};
		rom[ 732  ] = { 5'd16,	5'd12,	5'd6,	5'd4};
		rom[ 733  ] = { 5'd2,	5'd12,	5'd6,	5'd4};
		rom[ 734  ] = { 5'd10,	5'd7,	5'd4,	5'd5};
		rom[ 735  ] = { 5'd1,	5'd6,	5'd19,	5'd1};
		rom[ 736  ] = { 5'd14,	5'd8,	5'd3,	5'd7};
		rom[ 737  ] = { 5'd3,	5'd11,	5'd12,	5'd3};
		rom[ 738  ] = { 5'd3,	5'd7,	5'd18,	5'd1};
		rom[ 739  ] = { 5'd10,	5'd6,	5'd4,	5'd6};
		rom[ 740  ] = { 5'd3,	5'd9,	5'd9,	5'd14};
		rom[ 741  ] = { 5'd2,	5'd0,	5'd2,	5'd9};
		rom[ 742  ] = { 5'd12,	5'd5,	5'd2,	5'd18};
		rom[ 743  ] = { 5'd10,	5'd5,	5'd2,	5'd18};
		rom[ 744  ] = { 5'd12,	5'd5,	5'd2,	5'd10};
		rom[ 745  ] = { 5'd11,	5'd4,	5'd2,	5'd11};
		rom[ 746  ] = { 5'd4,	5'd17,	5'd18,	5'd1};
		rom[ 747  ] = { 5'd0,	5'd17,	5'd20,	5'd1};
		rom[ 748  ] = { 5'd9,	5'd13,	5'd6,	5'd4};
		rom[ 749  ] = { 5'd8,	5'd17,	5'd8,	5'd4};
		rom[ 750  ] = { 5'd13,	5'd16,	5'd3,	5'd6};
		rom[ 751  ] = { 5'd5,	5'd9,	5'd7,	5'd7};
		rom[ 752  ] = { 5'd12,	5'd0,	5'd12,	5'd5};
		rom[ 753  ] = { 5'd1,	5'd12,	5'd18,	5'd1};
		rom[ 754  ] = { 5'd19,	5'd9,	5'd5,	5'd4};
		rom[ 755  ] = { 5'd0,	5'd9,	5'd5,	5'd4};
		rom[ 756  ] = { 5'd20,	5'd6,	5'd4,	5'd9};
		rom[ 757  ] = { 5'd0,	5'd6,	5'd4,	5'd9};
		rom[ 758  ] = { 5'd18,	5'd5,	5'd6,	5'd6};
		rom[ 759  ] = { 5'd9,	5'd6,	5'd2,	5'd9};
		rom[ 760  ] = { 5'd11,	5'd13,	5'd2,	5'd11};
		rom[ 761  ] = { 5'd0,	5'd5,	5'd6,	5'd6};
		rom[ 762  ] = { 5'd1,	5'd3,	5'd23,	5'd1};
		rom[ 763  ] = { 5'd1,	5'd16,	5'd19,	5'd1};
		rom[ 764  ] = { 5'd13,	5'd19,	5'd11,	5'd2};
		rom[ 765  ] = { 5'd4,	5'd13,	5'd4,	5'd5};
		rom[ 766  ] = { 5'd12,	5'd10,	5'd5,	5'd4};
		rom[ 767  ] = { 5'd4,	5'd9,	5'd9,	5'd3};
		rom[ 768  ] = { 5'd15,	5'd16,	5'd9,	5'd2};
		rom[ 769  ] = { 5'd1,	5'd14,	5'd9,	5'd2};
		rom[ 770  ] = { 5'd13,	5'd10,	5'd10,	5'd4};
		rom[ 771  ] = { 5'd5,	5'd0,	5'd3,	5'd18};
		rom[ 772  ] = { 5'd16,	5'd11,	5'd3,	5'd10};
		rom[ 773  ] = { 5'd5,	5'd2,	5'd4,	5'd5};
		rom[ 774  ] = { 5'd10,	5'd4,	5'd7,	5'd6};
		rom[ 775  ] = { 5'd7,	5'd0,	5'd5,	5'd7};
		rom[ 776  ] = { 5'd12,	5'd19,	5'd12,	5'd2};
		rom[ 777  ] = { 5'd0,	5'd8,	5'd23,	5'd2};
		rom[ 778  ] = { 5'd17,	5'd10,	5'd4,	5'd5};
		rom[ 779  ] = { 5'd0,	5'd17,	5'd18,	5'd1};
		rom[ 780  ] = { 5'd15,	5'd18,	5'd9,	5'd2};
		rom[ 781  ] = { 5'd0,	5'd18,	5'd9,	5'd2};
		rom[ 782  ] = { 5'd13,	5'd11,	5'd3,	5'd6};
		rom[ 783  ] = { 5'd8,	5'd11,	5'd3,	5'd6};
		rom[ 784  ] = { 5'd12,	5'd3,	5'd12,	5'd3};
		rom[ 785  ] = { 5'd2,	5'd5,	5'd18,	5'd1};
		rom[ 786  ] = { 5'd12,	5'd0,	5'd12,	5'd2};
		rom[ 787  ] = { 5'd1,	5'd17,	5'd18,	5'd1};
		rom[ 788  ] = { 5'd15,	5'd17,	5'd9,	5'd2};
		rom[ 789  ] = { 5'd0,	5'd17,	5'd9,	5'd2};
		rom[ 790  ] = { 5'd6,	5'd18,	5'd18,	5'd1};
		rom[ 791  ] = { 5'd10,	5'd8,	5'd2,	5'd10};
		rom[ 792  ] = { 5'd12,	5'd6,	5'd2,	5'd9};
		rom[ 793  ] = { 5'd8,	5'd12,	5'd5,	5'd4};
		rom[ 794  ] = { 5'd12,	5'd12,	5'd6,	5'd4};
		rom[ 795  ] = { 5'd8,	5'd5,	5'd2,	5'd11};
		rom[ 796  ] = { 5'd13,	5'd9,	5'd8,	5'd3};
		rom[ 797  ] = { 5'd1,	5'd9,	5'd21,	5'd2};
		rom[ 798  ] = { 5'd15,	5'd11,	5'd3,	5'd6};
		rom[ 799  ] = { 5'd6,	5'd13,	5'd11,	5'd4};
		rom[ 800  ] = { 5'd18,	5'd8,	5'd5,	5'd4};
		rom[ 801  ] = { 5'd11,	5'd8,	5'd6,	5'd3};
		rom[ 802  ] = { 5'd12,	5'd11,	5'd6,	5'd4};
		rom[ 803  ] = { 5'd0,	5'd11,	5'd22,	5'd11};
		rom[ 804  ] = { 5'd11,	5'd6,	5'd6,	5'd4};
		rom[ 805  ] = { 5'd11,	5'd0,	5'd2,	5'd9};
		rom[ 806  ] = { 5'd12,	5'd0,	5'd2,	5'd9};
		rom[ 807  ] = { 5'd8,	5'd3,	5'd3,	5'd7};
		rom[ 808  ] = { 5'd9,	5'd10,	5'd6,	5'd8};
		rom[ 809  ] = { 5'd10,	5'd7,	5'd3,	5'd7};
		rom[ 810  ] = { 5'd4,	5'd13,	5'd16,	5'd10};
		rom[ 811  ] = { 5'd11,	5'd4,	5'd2,	5'd10};
		rom[ 812  ] = { 5'd5,	5'd2,	5'd16,	5'd2};
		rom[ 813  ] = { 5'd8,	5'd5,	5'd6,	5'd4};
		rom[ 814  ] = { 5'd15,	5'd0,	5'd2,	5'd9};
		rom[ 815  ] = { 5'd12,	5'd4,	5'd4,	5'd5};
		rom[ 816  ] = { 5'd12,	5'd10,	5'd5,	5'd4};
		rom[ 817  ] = { 5'd7,	5'd10,	5'd5,	5'd4};
		rom[ 818  ] = { 5'd11,	5'd11,	5'd4,	5'd5};
		rom[ 819  ] = { 5'd3,	5'd10,	5'd4,	5'd5};
		rom[ 820  ] = { 5'd14,	5'd12,	5'd3,	5'd8};
		rom[ 821  ] = { 5'd8,	5'd21,	5'd8,	5'd3};
		rom[ 822  ] = { 5'd9,	5'd20,	5'd6,	5'd4};
		rom[ 823  ] = { 5'd1,	5'd17,	5'd9,	5'd2};
		rom[ 824  ] = { 5'd11,	5'd19,	5'd10,	5'd2};
		rom[ 825  ] = { 5'd9,	5'd18,	5'd4,	5'd6};
		rom[ 826  ] = { 5'd12,	5'd6,	5'd3,	5'd6};
		rom[ 827  ] = { 5'd1,	5'd16,	5'd6,	5'd3};
		rom[ 828  ] = { 5'd6,	5'd18,	5'd12,	5'd2};
		rom[ 829  ] = { 5'd1,	5'd6,	5'd20,	5'd1};
		rom[ 830  ] = { 5'd8,	5'd4,	5'd9,	5'd3};
		rom[ 831  ] = { 5'd2,	5'd21,	5'd9,	5'd2};
		rom[ 832  ] = { 5'd11,	5'd7,	5'd4,	5'd6};
		rom[ 833  ] = { 5'd7,	5'd2,	5'd4,	5'd6};
		rom[ 834  ] = { 5'd14,	5'd10,	5'd3,	5'd8};
		rom[ 835  ] = { 5'd9,	5'd11,	5'd4,	5'd5};
		rom[ 836  ] = { 5'd14,	5'd9,	5'd3,	5'd6};
		rom[ 837  ] = { 5'd7,	5'd10,	5'd2,	5'd9};
		rom[ 838  ] = { 5'd4,	5'd11,	5'd5,	5'd4};
		rom[ 839  ] = { 5'd9,	5'd0,	5'd7,	5'd6};
		rom[ 840  ] = { 5'd7,	5'd8,	5'd10,	5'd2};
		rom[ 841  ] = { 5'd11,	5'd0,	5'd2,	5'd15};
		rom[ 842  ] = { 5'd2,	5'd3,	5'd18,	5'd1};
		rom[ 843  ] = { 5'd8,	5'd20,	5'd8,	5'd3};
		rom[ 844  ] = { 5'd3,	5'd1,	5'd18,	5'd1};
		rom[ 845  ] = { 5'd11,	5'd0,	5'd3,	5'd6};
		rom[ 846  ] = { 5'd0,	5'd18,	5'd18,	5'd1};
		rom[ 847  ] = { 5'd10,	5'd7,	5'd4,	5'd5};
		rom[ 848  ] = { 5'd2,	5'd3,	5'd2,	5'd9};
		rom[ 849  ] = { 5'd20,	5'd2,	5'd2,	5'd9};
		rom[ 850  ] = { 5'd2,	5'd2,	5'd2,	5'd9};
		rom[ 851  ] = { 5'd12,	5'd1,	5'd12,	5'd2};
		rom[ 852  ] = { 5'd0,	5'd18,	5'd9,	5'd2};
		rom[ 853  ] = { 5'd14,	5'd15,	5'd9,	5'd2};
		rom[ 854  ] = { 5'd0,	5'd16,	5'd19,	5'd1};
		rom[ 855  ] = { 5'd12,	5'd5,	5'd11,	5'd6};
		rom[ 856  ] = { 5'd8,	5'd13,	5'd3,	5'd6};
		rom[ 857  ] = { 5'd4,	5'd3,	5'd20,	5'd1};
		rom[ 858  ] = { 5'd10,	5'd14,	5'd2,	5'd10};
		rom[ 859  ] = { 5'd14,	5'd12,	5'd8,	5'd3};
		rom[ 860  ] = { 5'd2,	5'd16,	5'd8,	5'd3};
		rom[ 861  ] = { 5'd14,	5'd8,	5'd3,	5'd7};
		rom[ 862  ] = { 5'd2,	5'd12,	5'd8,	5'd3};
		rom[ 863  ] = { 5'd5,	5'd20,	5'd16,	5'd4};
		rom[ 864  ] = { 5'd9,	5'd7,	5'd4,	5'd6};
		rom[ 865  ] = { 5'd12,	5'd2,	5'd4,	5'd5};
		rom[ 866  ] = { 5'd6,	5'd6,	5'd6,	5'd3};
		rom[ 867  ] = { 5'd12,	5'd7,	5'd2,	5'd9};
		rom[ 868  ] = { 5'd0,	5'd0,	5'd4,	5'd6};
		rom[ 869  ] = { 5'd18,	5'd11,	5'd6,	5'd3};
		rom[ 870  ] = { 5'd5,	5'd12,	5'd3,	5'd6};
		rom[ 871  ] = { 5'd10,	5'd21,	5'd7,	5'd3};
		rom[ 872  ] = { 5'd2,	5'd3,	5'd16,	5'd3};
		rom[ 873  ] = { 5'd13,	5'd9,	5'd7,	5'd3};
		rom[ 874  ] = { 5'd6,	5'd11,	5'd4,	5'd7};
		rom[ 875  ] = { 5'd11,	5'd7,	5'd2,	5'd9};
		rom[ 876  ] = { 5'd7,	5'd8,	5'd3,	5'd7};
		rom[ 877  ] = { 5'd18,	5'd16,	5'd4,	5'd8};
		rom[ 878  ] = { 5'd11,	5'd14,	5'd2,	5'd10};
		rom[ 879  ] = { 5'd10,	5'd11,	5'd4,	5'd5};
		rom[ 880  ] = { 5'd0,	5'd13,	5'd23,	5'd1};
		rom[ 881  ] = { 5'd15,	5'd0,	5'd2,	5'd12};
		rom[ 882  ] = { 5'd4,	5'd10,	5'd4,	5'd5};
		rom[ 883  ] = { 5'd13,	5'd4,	5'd10,	5'd2};
		rom[ 884  ] = { 5'd7,	5'd0,	5'd2,	5'd12};
		rom[ 885  ] = { 5'd14,	5'd6,	5'd3,	5'd6};
		rom[ 886  ] = { 5'd7,	5'd6,	5'd3,	5'd6};
		rom[ 887  ] = { 5'd12,	5'd11,	5'd6,	5'd13};
		rom[ 888  ] = { 5'd6,	5'd11,	5'd6,	5'd13};
		rom[ 889  ] = { 5'd16,	5'd16,	5'd4,	5'd6};
		rom[ 890  ] = { 5'd0,	5'd7,	5'd21,	5'd1};
		rom[ 891  ] = { 5'd16,	5'd16,	5'd4,	5'd6};
		rom[ 892  ] = { 5'd5,	5'd14,	5'd6,	5'd7};
		rom[ 893  ] = { 5'd5,	5'd11,	5'd19,	5'd1};
		rom[ 894  ] = { 5'd5,	5'd6,	5'd14,	5'd2};
		rom[ 895  ] = { 5'd9,	5'd18,	5'd6,	5'd4};
		rom[ 896  ] = { 5'd9,	5'd0,	5'd2,	5'd9};
		rom[ 897  ] = { 5'd13,	5'd5,	5'd11,	5'd2};
		rom[ 898  ] = { 5'd5,	5'd0,	5'd3,	5'd6};
		rom[ 899  ] = { 5'd19,	5'd1,	5'd2,	5'd23};
		rom[ 900  ] = { 5'd3,	5'd1,	5'd2,	5'd23};
		rom[ 901  ] = { 5'd5,	5'd17,	5'd18,	5'd1};
		rom[ 902  ] = { 5'd0,	5'd5,	5'd11,	5'd2};
		rom[ 903  ] = { 5'd2,	5'd17,	5'd20,	5'd1};
		rom[ 904  ] = { 5'd5,	5'd5,	5'd13,	5'd2};
		rom[ 905  ] = { 5'd1,	5'd9,	5'd11,	5'd15};
		rom[ 906  ] = { 5'd10,	5'd4,	5'd7,	5'd3};
		rom[ 907  ] = { 5'd8,	5'd7,	5'd5,	5'd4};
		rom[ 908  ] = { 5'd11,	5'd7,	5'd5,	5'd4};
		rom[ 909  ] = { 5'd12,	5'd4,	5'd2,	5'd9};
		rom[ 910  ] = { 5'd4,	5'd12,	5'd3,	5'd6};
		rom[ 911  ] = { 5'd12,	5'd3,	5'd4,	5'd5};
		rom[ 912  ] = { 5'd3,	5'd6,	5'd8,	5'd3};
		rom[ 913  ] = { 5'd5,	5'd9,	5'd14,	5'd3};
		rom[ 914  ] = { 5'd4,	5'd5,	5'd9,	5'd2};
		rom[ 915  ] = { 5'd6,	5'd4,	5'd18,	5'd1};
		rom[ 916  ] = { 5'd10,	5'd6,	5'd3,	5'd6};
		rom[ 917  ] = { 5'd0,	5'd2,	5'd24,	5'd1};
		rom[ 918  ] = { 5'd0,	5'd19,	5'd10,	5'd2};
		rom[ 919  ] = { 5'd3,	5'd19,	5'd18,	5'd1};
		rom[ 920  ] = { 5'd2,	5'd5,	5'd3,	5'd8};
		rom[ 921  ] = { 5'd7,	5'd8,	5'd11,	5'd2};
		rom[ 922  ] = { 5'd5,	5'd13,	5'd12,	5'd11};
		rom[ 923  ] = { 5'd10,	5'd12,	5'd4,	5'd5};
		rom[ 924  ] = { 5'd9,	5'd6,	5'd4,	5'd6};
		rom[ 925  ] = { 5'd18,	5'd11,	5'd6,	5'd3};
		rom[ 926  ] = { 5'd9,	5'd7,	5'd5,	5'd10};
		rom[ 927  ] = { 5'd12,	5'd5,	5'd2,	5'd9};
		rom[ 928  ] = { 5'd11,	5'd9,	5'd2,	5'd10};
		rom[ 929  ] = { 5'd13,	5'd14,	5'd2,	5'd10};
		rom[ 930  ] = { 5'd9,	5'd14,	5'd2,	5'd10};
		rom[ 931  ] = { 5'd4,	5'd11,	5'd16,	5'd3};
		rom[ 932  ] = { 5'd2,	5'd12,	5'd20,	5'd1};
		rom[ 933  ] = { 5'd13,	5'd0,	5'd2,	5'd13};
		rom[ 934  ] = { 5'd9,	5'd0,	5'd2,	5'd13};
		rom[ 935  ] = { 5'd9,	5'd1,	5'd6,	5'd7};
		rom[ 936  ] = { 5'd1,	5'd14,	5'd6,	5'd3};
		rom[ 937  ] = { 5'd8,	5'd20,	5'd9,	5'd2};
		rom[ 938  ] = { 5'd3,	5'd11,	5'd15,	5'd2};
		rom[ 939  ] = { 5'd5,	5'd11,	5'd19,	5'd1};
		rom[ 940  ] = { 5'd8,	5'd14,	5'd7,	5'd8};
		rom[ 941  ] = { 5'd9,	5'd16,	5'd9,	5'd2};
		rom[ 942  ] = { 5'd0,	5'd11,	5'd8,	5'd4};
		rom[ 943  ] = { 5'd6,	5'd5,	5'd18,	5'd1};
		rom[ 944  ] = { 5'd4,	5'd16,	5'd4,	5'd6};
		rom[ 945  ] = { 5'd13,	5'd15,	5'd9,	5'd2};
		rom[ 946  ] = { 5'd5,	5'd8,	5'd7,	5'd7};
		rom[ 947  ] = { 5'd12,	5'd16,	5'd11,	5'd3};
		rom[ 948  ] = { 5'd11,	5'd0,	5'd2,	5'd9};
		rom[ 949  ] = { 5'd14,	5'd5,	5'd5,	5'd5};
		rom[ 950  ] = { 5'd5,	5'd5,	5'd5,	5'd5};
		rom[ 951  ] = { 5'd12,	5'd6,	5'd8,	5'd3};
		rom[ 952  ] = { 5'd0,	5'd10,	5'd6,	5'd3};
		rom[ 953  ] = { 5'd20,	5'd10,	5'd4,	5'd7};
		rom[ 954  ] = { 5'd9,	5'd18,	5'd6,	5'd6};
		rom[ 955  ] = { 5'd12,	5'd10,	5'd4,	5'd6};
		rom[ 956  ] = { 5'd10,	5'd0,	5'd2,	5'd9};
		rom[ 957  ] = { 5'd14,	5'd4,	5'd4,	5'd8};
		rom[ 958  ] = { 5'd7,	5'd12,	5'd10,	5'd2};
		rom[ 959  ] = { 5'd12,	5'd6,	5'd7,	5'd7};
		rom[ 960  ] = { 5'd2,	5'd12,	5'd20,	5'd1};
		rom[ 961  ] = { 5'd18,	5'd16,	5'd4,	5'd8};
		rom[ 962  ] = { 5'd1,	5'd11,	5'd6,	5'd5};
		rom[ 963  ] = { 5'd6,	5'd11,	5'd12,	5'd2};
		rom[ 964  ] = { 5'd12,	5'd12,	5'd3,	5'd7};
		rom[ 965  ] = { 5'd14,	5'd4,	5'd4,	5'd8};
		rom[ 966  ] = { 5'd6,	5'd4,	5'd4,	5'd8};
		rom[ 967  ] = { 5'd11,	5'd9,	5'd3,	5'd6};
		rom[ 968  ] = { 5'd1,	5'd5,	5'd8,	5'd6};
		rom[ 969  ] = { 5'd9,	5'd9,	5'd3,	5'd8};
		rom[ 970  ] = { 5'd7,	5'd0,	5'd1,	5'd18};
		rom[ 971  ] = { 5'd17,	5'd16,	5'd5,	5'd7};
		rom[ 972  ] = { 5'd2,	5'd16,	5'd5,	5'd7};
		rom[ 973  ] = { 5'd7,	5'd7,	5'd10,	5'd3};
		rom[ 974  ] = { 5'd1,	5'd9,	5'd23,	5'd6};
		rom[ 975  ] = { 5'd8,	5'd1,	5'd7,	5'd3};
		rom[ 976  ] = { 5'd11,	5'd6,	5'd2,	5'd9};
		rom[ 977  ] = { 5'd3,	5'd18,	5'd6,	5'd3};
		rom[ 978  ] = { 5'd20,	5'd8,	5'd4,	5'd8};
		rom[ 979  ] = { 5'd8,	5'd19,	5'd8,	5'd4};
		rom[ 980  ] = { 5'd20,	5'd8,	5'd4,	5'd8};
		rom[ 981  ] = { 5'd0,	5'd8,	5'd4,	5'd8};
		rom[ 982  ] = { 5'd8,	5'd17,	5'd8,	5'd5};
		rom[ 983  ] = { 5'd5,	5'd11,	5'd5,	5'd4};
		rom[ 984  ] = { 5'd4,	5'd2,	5'd19,	5'd1};
		rom[ 985  ] = { 5'd8,	5'd12,	5'd8,	5'd9};
		rom[ 986  ] = { 5'd6,	5'd4,	5'd13,	5'd4};
		rom[ 987  ] = { 5'd0,	5'd1,	5'd24,	5'd1};
		rom[ 988  ] = { 5'd20,	5'd3,	5'd2,	5'd11};
		rom[ 989  ] = { 5'd10,	5'd6,	5'd2,	5'd9};
		rom[ 990  ] = { 5'd12,	5'd11,	5'd6,	5'd4};
		rom[ 991  ] = { 5'd0,	5'd8,	5'd6,	5'd3};
		rom[ 992  ] = { 5'd6,	5'd18,	5'd18,	5'd1};
		rom[ 993  ] = { 5'd0,	5'd16,	5'd9,	5'd2};
		rom[ 994  ] = { 5'd20,	5'd3,	5'd2,	5'd9};
		rom[ 995  ] = { 5'd2,	5'd3,	5'd2,	5'd9};
		rom[ 996  ] = { 5'd18,	5'd0,	5'd3,	5'd19};
		rom[ 997  ] = { 5'd3,	5'd0,	5'd3,	5'd19};
		rom[ 998  ] = { 5'd13,	5'd11,	5'd3,	5'd8};
		rom[ 999  ] = { 5'd8,	5'd11,	5'd3,	5'd8};
		rom[ 1000 ] = { 5'd5,	5'd12,	5'd19,	5'd1};
		rom[ 1001 ] = { 5'd9,	5'd20,	5'd6,	5'd4};
		rom[ 1002 ] = { 5'd6,	5'd8,	5'd16,	5'd2};
		rom[ 1003 ] = { 5'd9,	5'd0,	5'd3,	5'd6};
		rom[ 1004 ] = { 5'd10,	5'd10,	5'd4,	5'd7};
		rom[ 1005 ] = { 5'd1,	5'd11,	5'd15,	5'd6};
		rom[ 1006 ] = { 5'd11,	5'd12,	5'd4,	5'd5};
		rom[ 1007 ] = { 5'd7,	5'd0,	5'd2,	5'd9};
		rom[ 1008 ] = { 5'd14,	5'd0,	5'd2,	5'd9};
		rom[ 1009 ] = { 5'd5,	5'd5,	5'd6,	5'd4};
		rom[ 1010 ] = { 5'd13,	5'd14,	5'd11,	5'd2};
		rom[ 1011 ] = { 5'd0,	5'd14,	5'd21,	5'd1};
		rom[ 1012 ] = { 5'd12,	5'd1,	5'd4,	5'd6};
		rom[ 1013 ] = { 5'd1,	5'd0,	5'd3,	5'd6};
		rom[ 1014 ] = { 5'd2,	5'd3,	5'd21,	5'd1};
		rom[ 1015 ] = { 5'd2,	5'd3,	5'd19,	5'd1};
		rom[ 1016 ] = { 5'd20,	5'd10,	5'd3,	5'd7};
		rom[ 1017 ] = { 5'd1,	5'd10,	5'd3,	5'd7};
		rom[ 1018 ] = { 5'd14,	5'd6,	5'd7,	5'd7};
		rom[ 1019 ] = { 5'd0,	5'd14,	5'd9,	5'd2};
		rom[ 1020 ] = { 5'd15,	5'd17,	5'd8,	5'd3};
		rom[ 1021 ] = { 5'd1,	5'd1,	5'd11,	5'd2};
		rom[ 1022 ] = { 5'd9,	5'd13,	5'd9,	5'd2};
		rom[ 1023 ] = { 5'd0,	5'd16,	5'd18,	5'd1};
		rom[ 1024 ] = { 5'd16,	5'd17,	5'd7,	5'd3};
		rom[ 1025 ] = { 5'd12,	5'd3,	5'd8,	5'd4};
		rom[ 1026 ] = { 5'd7,	5'd6,	5'd6,	5'd5};
		rom[ 1027 ] = { 5'd11,	5'd6,	5'd2,	5'd9};
		rom[ 1028 ] = { 5'd12,	5'd1,	5'd2,	5'd10};
		rom[ 1029 ] = { 5'd10,	5'd1,	5'd2,	5'd10};
		rom[ 1030 ] = { 5'd15,	5'd18,	5'd6,	5'd3};
		rom[ 1031 ] = { 5'd3,	5'd18,	5'd6,	5'd3};
		rom[ 1032 ] = { 5'd16,	5'd1,	5'd1,	5'd19};
		rom[ 1033 ] = { 5'd3,	5'd3,	5'd2,	5'd9};
		rom[ 1034 ] = { 5'd16,	5'd0,	5'd1,	5'd19};
		rom[ 1035 ] = { 5'd12,	5'd3,	5'd6,	5'd4};
		rom[ 1036 ] = { 5'd10,	5'd5,	5'd2,	5'd9};
		rom[ 1037 ] = { 5'd7,	5'd0,	5'd1,	5'd19};
		rom[ 1038 ] = { 5'd11,	5'd7,	5'd3,	5'd6};
		rom[ 1039 ] = { 5'd11,	5'd7,	5'd5,	5'd5};
		rom[ 1040 ] = { 5'd12,	5'd3,	5'd1,	5'd18};
		rom[ 1041 ] = { 5'd11,	5'd3,	5'd2,	5'd12};
		rom[ 1042 ] = { 5'd3,	5'd8,	5'd19,	5'd1};
		rom[ 1043 ] = { 5'd2,	5'd8,	5'd18,	5'd1};
		rom[ 1044 ] = { 5'd12,	5'd13,	5'd9,	5'd2};
		rom[ 1045 ] = { 5'd5,	5'd5,	5'd2,	5'd9};
		rom[ 1046 ] = { 5'd14,	5'd1,	5'd10,	5'd2};
		rom[ 1047 ] = { 5'd0,	5'd1,	5'd10,	5'd2};
		rom[ 1048 ] = { 5'd10,	5'd15,	5'd3,	5'd6};
		rom[ 1049 ] = { 5'd8,	5'd2,	5'd8,	5'd8};
		rom[ 1050 ] = { 5'd5,	5'd6,	5'd18,	5'd1};
		rom[ 1051 ] = { 5'd11,	5'd15,	5'd3,	5'd6};
		rom[ 1052 ] = { 5'd11,	5'd12,	5'd4,	5'd5};
		rom[ 1053 ] = { 5'd9,	5'd12,	5'd4,	5'd5};
		rom[ 1054 ] = { 5'd5,	5'd2,	5'd14,	5'd2};
		rom[ 1055 ] = { 5'd10,	5'd7,	5'd4,	5'd5};
		rom[ 1056 ] = { 5'd10,	5'd11,	5'd5,	5'd4};
		rom[ 1057 ] = { 5'd7,	5'd9,	5'd4,	5'd7};
		rom[ 1058 ] = { 5'd12,	5'd5,	5'd11,	5'd3};
		rom[ 1059 ] = { 5'd0,	5'd8,	5'd6,	5'd3};
		rom[ 1060 ] = { 5'd12,	5'd19,	5'd9,	5'd2};
		rom[ 1061 ] = { 5'd2,	5'd19,	5'd19,	5'd1};
		rom[ 1062 ] = { 5'd12,	5'd19,	5'd9,	5'd2};
		rom[ 1063 ] = { 5'd1,	5'd18,	5'd18,	5'd1};
		rom[ 1064 ] = { 5'd12,	5'd19,	5'd9,	5'd2};
		rom[ 1065 ] = { 5'd0,	5'd1,	5'd24,	5'd1};
		rom[ 1066 ] = { 5'd5,	5'd2,	5'd14,	5'd2};
		rom[ 1067 ] = { 5'd6,	5'd16,	5'd9,	5'd2};
		rom[ 1068 ] = { 5'd14,	5'd16,	5'd6,	5'd3};
		rom[ 1069 ] = { 5'd5,	5'd22,	5'd13,	5'd2};
		rom[ 1070 ] = { 5'd9,	5'd13,	5'd6,	5'd4};
		rom[ 1071 ] = { 5'd8,	5'd10,	5'd7,	5'd3};
		rom[ 1072 ] = { 5'd11,	5'd8,	5'd3,	5'd6};
		rom[ 1073 ] = { 5'd6,	5'd10,	5'd3,	5'd7};
		rom[ 1074 ] = { 5'd17,	5'd10,	5'd5,	5'd4};
		rom[ 1075 ] = { 5'd8,	5'd15,	5'd8,	5'd3};
		rom[ 1076 ] = { 5'd8,	5'd7,	5'd9,	5'd2};
		rom[ 1077 ] = { 5'd4,	5'd16,	5'd6,	5'd3};
		rom[ 1078 ] = { 5'd12,	5'd19,	5'd9,	5'd2};
		rom[ 1079 ] = { 5'd9,	5'd15,	5'd6,	5'd3};
		rom[ 1080 ] = { 5'd16,	5'd9,	5'd7,	5'd5};
		rom[ 1081 ] = { 5'd1,	5'd9,	5'd7,	5'd5};
		rom[ 1082 ] = { 5'd11,	5'd7,	5'd3,	5'd17};
		rom[ 1083 ] = { 5'd3,	5'd4,	5'd3,	5'd10};
		rom[ 1084 ] = { 5'd7,	5'd8,	5'd5,	5'd4};
		rom[ 1085 ] = { 5'd12,	5'd7,	5'd2,	5'd9};
		rom[ 1086 ] = { 5'd12,	5'd15,	5'd2,	5'd9};
		rom[ 1087 ] = { 5'd3,	5'd8,	5'd3,	5'd8};
		rom[ 1088 ] = { 5'd12,	5'd19,	5'd9,	5'd2};
		rom[ 1089 ] = { 5'd3,	5'd19,	5'd9,	5'd2};
		rom[ 1090 ] = { 5'd13,	5'd1,	5'd3,	5'd6};
		rom[ 1091 ] = { 5'd5,	5'd12,	5'd4,	5'd5};
		rom[ 1092 ] = { 5'd11,	5'd5,	5'd4,	5'd6};
		rom[ 1093 ] = { 5'd9,	5'd4,	5'd3,	5'd8};
		rom[ 1094 ] = { 5'd17,	5'd16,	5'd5,	5'd4};
		rom[ 1095 ] = { 5'd2,	5'd16,	5'd5,	5'd4};
		rom[ 1096 ] = { 5'd12,	5'd0,	5'd12,	5'd2};
		rom[ 1097 ] = { 5'd0,	5'd8,	5'd9,	5'd2};
		rom[ 1098 ] = { 5'd12,	5'd4,	5'd12,	5'd3};
		rom[ 1099 ] = { 5'd5,	5'd2,	5'd11,	5'd2};
		rom[ 1100 ] = { 5'd12,	5'd1,	5'd11,	5'd2};
		rom[ 1101 ] = { 5'd9,	5'd15,	5'd6,	5'd9};
		rom[ 1102 ] = { 5'd2,	5'd11,	5'd20,	5'd2};
		rom[ 1103 ] = { 5'd5,	5'd9,	5'd14,	5'd7};
		rom[ 1104 ] = { 5'd4,	5'd5,	5'd16,	5'd3};
		rom[ 1105 ] = { 5'd2,	5'd4,	5'd19,	5'd1};
		rom[ 1106 ] = { 5'd7,	5'd3,	5'd10,	5'd2};
		rom[ 1107 ] = { 5'd0,	5'd14,	5'd4,	5'd5};
		rom[ 1108 ] = { 5'd2,	5'd11,	5'd21,	5'd1};
		rom[ 1109 ] = { 5'd6,	5'd0,	5'd3,	5'd6};
		rom[ 1110 ] = { 5'd6,	5'd7,	5'd14,	5'd3};
		rom[ 1111 ] = { 5'd11,	5'd1,	5'd2,	5'd9};
		rom[ 1112 ] = { 5'd15,	5'd11,	5'd9,	5'd3};
		rom[ 1113 ] = { 5'd8,	5'd7,	5'd4,	5'd7};
		rom[ 1114 ] = { 5'd3,	5'd23,	5'd19,	5'd1};
		rom[ 1115 ] = { 5'd2,	5'd16,	5'd20,	5'd1};
		rom[ 1116 ] = { 5'd19,	5'd0,	5'd2,	5'd13};
		rom[ 1117 ] = { 5'd1,	5'd11,	5'd8,	5'd4};
		rom[ 1118 ] = { 5'd14,	5'd17,	5'd6,	5'd3};
		rom[ 1119 ] = { 5'd4,	5'd17,	5'd6,	5'd3};
		rom[ 1120 ] = { 5'd14,	5'd5,	5'd2,	5'd10};
		rom[ 1121 ] = { 5'd8,	5'd5,	5'd2,	5'd10};
		rom[ 1122 ] = { 5'd14,	5'd8,	5'd6,	5'd3};
		rom[ 1123 ] = { 5'd4,	5'd8,	5'd6,	5'd3};
		rom[ 1124 ] = { 5'd8,	5'd2,	5'd8,	5'd21};
		rom[ 1125 ] = { 5'd3,	5'd2,	5'd2,	5'd13};
		rom[ 1126 ] = { 5'd20,	5'd0,	5'd2,	5'd21};
		rom[ 1127 ] = { 5'd2,	5'd4,	5'd2,	5'd20};
		rom[ 1128 ] = { 5'd8,	5'd18,	5'd9,	5'd2};
		rom[ 1129 ] = { 5'd9,	5'd0,	5'd2,	5'd9};
		rom[ 1130 ] = { 5'd16,	5'd15,	5'd7,	5'd3};
		rom[ 1131 ] = { 5'd12,	5'd21,	5'd7,	5'd3};
		rom[ 1132 ] = { 5'd11,	5'd5,	5'd3,	5'd9};
		rom[ 1133 ] = { 5'd12,	5'd5,	5'd2,	5'd10};
		rom[ 1134 ] = { 5'd12,	5'd6,	5'd2,	5'd9};
		rom[ 1135 ] = { 5'd10,	5'd5,	5'd3,	5'd9};
		rom[ 1136 ] = { 5'd14,	5'd16,	5'd10,	5'd2};
		rom[ 1137 ] = { 5'd5,	5'd5,	5'd7,	5'd7};
		rom[ 1138 ] = { 5'd18,	5'd8,	5'd6,	5'd3};
		rom[ 1139 ] = { 5'd6,	5'd6,	5'd6,	5'd6};
		rom[ 1140 ] = { 5'd13,	5'd13,	5'd2,	5'd10};
		rom[ 1141 ] = { 5'd1,	5'd10,	5'd10,	5'd4};
		rom[ 1142 ] = { 5'd15,	5'd15,	5'd9,	5'd2};
		rom[ 1143 ] = { 5'd9,	5'd3,	5'd6,	5'd3};
		rom[ 1144 ] = { 5'd10,	5'd8,	5'd5,	5'd7};
		rom[ 1145 ] = { 5'd3,	5'd6,	5'd16,	5'd2};
		rom[ 1146 ] = { 5'd16,	5'd6,	5'd8,	5'd3};
		rom[ 1147 ] = { 5'd9,	5'd13,	5'd2,	5'd10};
		rom[ 1148 ] = { 5'd15,	5'd15,	5'd9,	5'd2};
		rom[ 1149 ] = { 5'd0,	5'd15,	5'd9,	5'd2};
		rom[ 1150 ] = { 5'd13,	5'd18,	5'd9,	5'd2};
		rom[ 1151 ] = { 5'd2,	5'd18,	5'd9,	5'd2};
		rom[ 1152 ] = { 5'd5,	5'd17,	5'd18,	5'd1};
		rom[ 1153 ] = { 5'd1,	5'd17,	5'd18,	5'd1};
		rom[ 1154 ] = { 5'd5,	5'd1,	5'd18,	5'd1};
		rom[ 1155 ] = { 5'd1,	5'd2,	5'd19,	5'd1};
		rom[ 1156 ] = { 5'd16,	5'd2,	5'd2,	5'd11};
		rom[ 1157 ] = { 5'd9,	5'd15,	5'd5,	5'd6};
		rom[ 1158 ] = { 5'd16,	5'd2,	5'd2,	5'd11};
		rom[ 1159 ] = { 5'd6,	5'd2,	5'd2,	5'd11};
		rom[ 1160 ] = { 5'd18,	5'd5,	5'd6,	5'd3};
		rom[ 1161 ] = { 5'd1,	5'd2,	5'd11,	5'd2};
		rom[ 1162 ] = { 5'd9,	5'd0,	5'd7,	5'd12};
		rom[ 1163 ] = { 5'd0,	5'd13,	5'd18,	5'd1};
		rom[ 1164 ] = { 5'd14,	5'd2,	5'd2,	5'd9};
		rom[ 1165 ] = { 5'd3,	5'd11,	5'd18,	5'd1};
		rom[ 1166 ] = { 5'd16,	5'd6,	5'd8,	5'd3};
		rom[ 1167 ] = { 5'd3,	5'd8,	5'd18,	5'd1};
		rom[ 1168 ] = { 5'd11,	5'd11,	5'd2,	5'd9};
		rom[ 1169 ] = { 5'd11,	5'd8,	5'd2,	5'd9};
		rom[ 1170 ] = { 5'd15,	5'd0,	5'd1,	5'd18};
		rom[ 1171 ] = { 5'd8,	5'd0,	5'd1,	5'd18};
		rom[ 1172 ] = { 5'd17,	5'd6,	5'd7,	5'd3};
		rom[ 1173 ] = { 5'd3,	5'd20,	5'd9,	5'd2};
		rom[ 1174 ] = { 5'd3,	5'd19,	5'd21,	5'd1};
		rom[ 1175 ] = { 5'd0,	5'd6,	5'd7,	5'd3};
		rom[ 1176 ] = { 5'd2,	5'd8,	5'd22,	5'd1};
		rom[ 1177 ] = { 5'd0,	5'd3,	5'd12,	5'd8};
		rom[ 1178 ] = { 5'd13,	5'd19,	5'd9,	5'd2};
		rom[ 1179 ] = { 5'd5,	5'd5,	5'd6,	5'd4};
		rom[ 1180 ] = { 5'd12,	5'd6,	5'd7,	5'd3};
		rom[ 1181 ] = { 5'd5,	5'd16,	5'd7,	5'd3};
		rom[ 1182 ] = { 5'd18,	5'd5,	5'd6,	5'd3};
		rom[ 1183 ] = { 5'd0,	5'd5,	5'd6,	5'd3};
		rom[ 1184 ] = { 5'd13,	5'd4,	5'd10,	5'd5};
		rom[ 1185 ] = { 5'd5,	5'd13,	5'd3,	5'd8};
		rom[ 1186 ] = { 5'd9,	5'd1,	5'd7,	5'd15};
		rom[ 1187 ] = { 5'd12,	5'd12,	5'd7,	5'd8};
		rom[ 1188 ] = { 5'd6,	5'd7,	5'd6,	5'd4};
		rom[ 1189 ] = { 5'd9,	5'd5,	5'd3,	5'd6};
		rom[ 1190 ] = { 5'd13,	5'd11,	5'd3,	5'd6};
		rom[ 1191 ] = { 5'd8,	5'd11,	5'd3,	5'd6};
		rom[ 1192 ] = { 5'd6,	5'd5,	5'd18,	5'd1};
		rom[ 1193 ] = { 5'd2,	5'd2,	5'd2,	5'd11};
		rom[ 1194 ] = { 5'd20,	5'd0,	5'd2,	5'd15};
		rom[ 1195 ] = { 5'd2,	5'd0,	5'd2,	5'd13};
		rom[ 1196 ] = { 5'd14,	5'd0,	5'd2,	5'd9};
		rom[ 1197 ] = { 5'd8,	5'd0,	5'd2,	5'd9};
		rom[ 1198 ] = { 5'd8,	5'd2,	5'd8,	5'd4};
		rom[ 1199 ] = { 5'd12,	5'd13,	5'd9,	5'd4};
		rom[ 1200 ] = { 5'd9,	5'd7,	5'd5,	5'd4};
		rom[ 1201 ] = { 5'd11,	5'd8,	5'd6,	5'd3};
		rom[ 1202 ] = { 5'd4,	5'd15,	5'd19,	5'd1};
		rom[ 1203 ] = { 5'd10,	5'd10,	5'd4,	5'd10};
		rom[ 1204 ] = { 5'd8,	5'd17,	5'd9,	5'd2};
		rom[ 1205 ] = { 5'd7,	5'd9,	5'd5,	5'd4};
		rom[ 1206 ] = { 5'd12,	5'd4,	5'd4,	5'd7};
		rom[ 1207 ] = { 5'd0,	5'd13,	5'd6,	5'd3};
		rom[ 1208 ] = { 5'd18,	5'd8,	5'd6,	5'd3};
		rom[ 1209 ] = { 5'd0,	5'd18,	5'd8,	5'd3};
		rom[ 1210 ] = { 5'd16,	5'd18,	5'd7,	5'd3};
		rom[ 1211 ] = { 5'd1,	5'd20,	5'd10,	5'd2};
		rom[ 1212 ] = { 5'd12,	5'd8,	5'd10,	5'd3};
		rom[ 1213 ] = { 5'd9,	5'd8,	5'd2,	5'd9};
		rom[ 1214 ] = { 5'd12,	5'd5,	5'd4,	5'd8};
		rom[ 1215 ] = { 5'd8,	5'd5,	5'd4,	5'd8};
		rom[ 1216 ] = { 5'd12,	5'd6,	5'd2,	5'd9};
		rom[ 1217 ] = { 5'd4,	5'd0,	5'd2,	5'd16};
		rom[ 1218 ] = { 5'd15,	5'd8,	5'd6,	5'd4};
		rom[ 1219 ] = { 5'd3,	5'd8,	5'd6,	5'd4};
		rom[ 1220 ] = { 5'd15,	5'd14,	5'd9,	5'd2};
		rom[ 1221 ] = { 5'd4,	5'd11,	5'd15,	5'd11};
		rom[ 1222 ] = { 5'd15,	5'd14,	5'd9,	5'd2};
		rom[ 1223 ] = { 5'd0,	5'd14,	5'd9,	5'd2};
		rom[ 1224 ] = { 5'd15,	5'd17,	5'd9,	5'd2};
		rom[ 1225 ] = { 5'd0,	5'd17,	5'd9,	5'd2};
		rom[ 1226 ] = { 5'd14,	5'd0,	5'd4,	5'd5};
		rom[ 1227 ] = { 5'd3,	5'd0,	5'd2,	5'd16};
		rom[ 1228 ] = { 5'd7,	5'd8,	5'd10,	5'd2};
		rom[ 1229 ] = { 5'd10,	5'd17,	5'd4,	5'd5};
		rom[ 1230 ] = { 5'd8,	5'd6,	5'd10,	5'd2};
		rom[ 1231 ] = { 5'd12,	5'd22,	5'd9,	5'd2};
		rom[ 1232 ] = { 5'd7,	5'd9,	5'd11,	5'd2};
		rom[ 1233 ] = { 5'd0,	5'd0,	5'd6,	5'd5};
		rom[ 1234 ] = { 5'd16,	5'd1,	5'd6,	5'd3};
		rom[ 1235 ] = { 5'd7,	5'd18,	5'd9,	5'd2};
		rom[ 1236 ] = { 5'd10,	5'd7,	5'd5,	5'd16};
		rom[ 1237 ] = { 5'd11,	5'd10,	5'd6,	5'd13};
		rom[ 1238 ] = { 5'd12,	5'd2,	5'd6,	5'd3};
		rom[ 1239 ] = { 5'd3,	5'd12,	5'd12,	5'd3};
		rom[ 1240 ] = { 5'd16,	5'd5,	5'd8,	5'd3};
		rom[ 1241 ] = { 5'd0,	5'd5,	5'd8,	5'd3};
		rom[ 1242 ] = { 5'd0,	5'd3,	5'd12,	5'd11};
		rom[ 1243 ] = { 5'd0,	5'd13,	5'd4,	5'd5};
		rom[ 1244 ] = { 5'd10,	5'd19,	5'd4,	5'd5};
		rom[ 1245 ] = { 5'd10,	5'd9,	5'd4,	5'd7};
		rom[ 1246 ] = { 5'd4,	5'd7,	5'd15,	5'd3};
		rom[ 1247 ] = { 5'd8,	5'd1,	5'd8,	5'd6};
		rom[ 1248 ] = { 5'd9,	5'd14,	5'd5,	5'd8};
		rom[ 1249 ] = { 5'd9,	5'd21,	5'd6,	5'd3};
		rom[ 1250 ] = { 5'd6,	5'd11,	5'd3,	5'd6};
		rom[ 1251 ] = { 5'd11,	5'd6,	5'd2,	5'd9};
		rom[ 1252 ] = { 5'd8,	5'd6,	5'd3,	5'd8};
		rom[ 1253 ] = { 5'd4,	5'd4,	5'd20,	5'd1};
		rom[ 1254 ] = { 5'd8,	5'd10,	5'd6,	5'd3};
		rom[ 1255 ] = { 5'd7,	5'd17,	5'd10,	5'd2};
		rom[ 1256 ] = { 5'd1,	5'd4,	5'd2,	5'd9};
		rom[ 1257 ] = { 5'd15,	5'd0,	5'd2,	5'd9};
		rom[ 1258 ] = { 5'd7,	5'd0,	5'd2,	5'd9};
		rom[ 1259 ] = { 5'd13,	5'd0,	5'd2,	5'd9};
		rom[ 1260 ] = { 5'd9,	5'd7,	5'd3,	5'd6};
		rom[ 1261 ] = { 5'd3,	5'd1,	5'd18,	5'd1};
		rom[ 1262 ] = { 5'd0,	5'd10,	5'd10,	5'd2};
		rom[ 1263 ] = { 5'd10,	5'd8,	5'd4,	5'd6};
		rom[ 1264 ] = { 5'd6,	5'd5,	5'd3,	5'd6};
		rom[ 1265 ] = { 5'd15,	5'd0,	5'd9,	5'd11};
		rom[ 1266 ] = { 5'd0,	5'd0,	5'd9,	5'd11};
		rom[ 1267 ] = { 5'd20,	5'd2,	5'd2,	5'd11};
		rom[ 1268 ] = { 5'd2,	5'd2,	5'd2,	5'd11};
		rom[ 1269 ] = { 5'd13,	5'd0,	5'd2,	5'd9};
		rom[ 1270 ] = { 5'd0,	5'd1,	5'd20,	5'd1};
		rom[ 1271 ] = { 5'd2,	5'd3,	5'd20,	5'd1};
		rom[ 1272 ] = { 5'd1,	5'd11,	5'd18,	5'd1};
		rom[ 1273 ] = { 5'd18,	5'd10,	5'd6,	5'd3};
		rom[ 1274 ] = { 5'd0,	5'd3,	5'd22,	5'd3};
		rom[ 1275 ] = { 5'd17,	5'd6,	5'd6,	5'd3};
		rom[ 1276 ] = { 5'd0,	5'd10,	5'd6,	5'd3};
		rom[ 1277 ] = { 5'd0,	5'd8,	5'd24,	5'd2};
		rom[ 1278 ] = { 5'd2,	5'd2,	5'd2,	5'd10};
		rom[ 1279 ] = { 5'd12,	5'd6,	5'd2,	5'd9};
		rom[ 1280 ] = { 5'd9,	5'd0,	5'd2,	5'd9};
		rom[ 1281 ] = { 5'd17,	5'd0,	5'd2,	5'd9};
		rom[ 1282 ] = { 5'd5,	5'd0,	5'd2,	5'd9};
		rom[ 1283 ] = { 5'd15,	5'd19,	5'd9,	5'd2};
		rom[ 1284 ] = { 5'd0,	5'd18,	5'd18,	5'd1};
		rom[ 1285 ] = { 5'd15,	5'd16,	5'd9,	5'd2};
		rom[ 1286 ] = { 5'd0,	5'd17,	5'd23,	5'd2};
		rom[ 1287 ] = { 5'd5,	5'd16,	5'd18,	5'd1};
		rom[ 1288 ] = { 5'd0,	5'd16,	5'd9,	5'd2};
		rom[ 1289 ] = { 5'd13,	5'd8,	5'd4,	5'd5};
		rom[ 1290 ] = { 5'd8,	5'd7,	5'd5,	5'd6};
		rom[ 1291 ] = { 5'd13,	5'd8,	5'd4,	5'd5};
		rom[ 1292 ] = { 5'd8,	5'd0,	5'd3,	5'd12};
		rom[ 1293 ] = { 5'd13,	5'd8,	5'd4,	5'd5};
		rom[ 1294 ] = { 5'd10,	5'd5,	5'd2,	5'd9};
		rom[ 1295 ] = { 5'd12,	5'd6,	5'd2,	5'd9};
		rom[ 1296 ] = { 5'd11,	5'd7,	5'd6,	5'd4};
		rom[ 1297 ] = { 5'd13,	5'd8,	5'd4,	5'd5};
		rom[ 1298 ] = { 5'd7,	5'd8,	5'd4,	5'd5};
		rom[ 1299 ] = { 5'd14,	5'd10,	5'd3,	5'd7};
		rom[ 1300 ] = { 5'd12,	5'd5,	5'd3,	5'd19};
		rom[ 1301 ] = { 5'd12,	5'd12,	5'd6,	5'd3};
		rom[ 1302 ] = { 5'd1,	5'd9,	5'd9,	5'd3};
		rom[ 1303 ] = { 5'd20,	5'd14,	5'd4,	5'd5};
		rom[ 1304 ] = { 5'd0,	5'd9,	5'd11,	5'd4};
		rom[ 1305 ] = { 5'd14,	5'd18,	5'd6,	5'd3};
		rom[ 1306 ] = { 5'd0,	5'd6,	5'd10,	5'd9};
		rom[ 1307 ] = { 5'd13,	5'd6,	5'd10,	5'd6};
		rom[ 1308 ] = { 5'd0,	5'd16,	5'd5,	5'd4};
		rom[ 1309 ] = { 5'd6,	5'd17,	5'd18,	5'd1};
		rom[ 1310 ] = { 5'd0,	5'd12,	5'd19,	5'd1};
		rom[ 1311 ] = { 5'd14,	5'd9,	5'd6,	5'd3};
		rom[ 1312 ] = { 5'd1,	5'd7,	5'd11,	5'd2};
		rom[ 1313 ] = { 5'd13,	5'd10,	5'd7,	5'd4};
		rom[ 1314 ] = { 5'd4,	5'd10,	5'd11,	5'd3};
		rom[ 1315 ] = { 5'd17,	5'd10,	5'd5,	5'd4};
		rom[ 1316 ] = { 5'd5,	5'd12,	5'd3,	5'd7};
		rom[ 1317 ] = { 5'd16,	5'd17,	5'd6,	5'd3};
		rom[ 1318 ] = { 5'd3,	5'd16,	5'd6,	5'd4};
		rom[ 1319 ] = { 5'd14,	5'd16,	5'd6,	5'd3};
		rom[ 1320 ] = { 5'd10,	5'd0,	5'd2,	5'd9};
		rom[ 1321 ] = { 5'd11,	5'd1,	5'd2,	5'd23};
		rom[ 1322 ] = { 5'd0,	5'd18,	5'd9,	5'd2};
		rom[ 1323 ] = { 5'd4,	5'd18,	5'd18,	5'd1};
		rom[ 1324 ] = { 5'd5,	5'd9,	5'd13,	5'd7};
		rom[ 1325 ] = { 5'd19,	5'd0,	5'd4,	5'd6};
		rom[ 1326 ] = { 5'd0,	5'd0,	5'd4,	5'd6};
		rom[ 1327 ] = { 5'd8,	5'd2,	5'd4,	5'd7};
		rom[ 1328 ] = { 5'd3,	5'd1,	5'd2,	5'd9};
		rom[ 1329 ] = { 5'd17,	5'd8,	5'd3,	5'd6};
		rom[ 1330 ] = { 5'd4,	5'd8,	5'd3,	5'd6};
		rom[ 1331 ] = { 5'd16,	5'd10,	5'd5,	5'd5};
		rom[ 1332 ] = { 5'd3,	5'd10,	5'd5,	5'd5};
		rom[ 1333 ] = { 5'd18,	5'd7,	5'd6,	5'd3};
		rom[ 1334 ] = { 5'd1,	5'd12,	5'd6,	5'd5};
		rom[ 1335 ] = { 5'd17,	5'd15,	5'd6,	5'd4};
		rom[ 1336 ] = { 5'd0,	5'd2,	5'd12,	5'd2};
		rom[ 1337 ] = { 5'd15,	5'd1,	5'd1,	5'd19};
		rom[ 1338 ] = { 5'd8,	5'd1,	5'd1,	5'd19};
		rom[ 1339 ] = { 5'd22,	5'd1,	5'd1,	5'd20};
		rom[ 1340 ] = { 5'd1,	5'd1,	5'd1,	5'd20};
		rom[ 1341 ] = { 5'd20,	5'd11,	5'd2,	5'd12};
		rom[ 1342 ] = { 5'd2,	5'd11,	5'd2,	5'd12};
		rom[ 1343 ] = { 5'd3,	5'd13,	5'd18,	5'd7};
		rom[ 1344 ] = { 5'd6,	5'd14,	5'd7,	5'd4};
		rom[ 1345 ] = { 5'd7,	5'd13,	5'd12,	5'd4};
		rom[ 1346 ] = { 5'd11,	5'd18,	5'd9,	5'd5};
		rom[ 1347 ] = { 5'd4,	5'd22,	5'd20,	5'd1};
		rom[ 1348 ] = { 5'd9,	5'd12,	5'd3,	5'd6};
		rom[ 1349 ] = { 5'd4,	5'd7,	5'd18,	5'd1};
		rom[ 1350 ] = { 5'd3,	5'd7,	5'd18,	5'd1};
		rom[ 1351 ] = { 5'd18,	5'd7,	5'd6,	5'd3};
		rom[ 1352 ] = { 5'd2,	5'd14,	5'd9,	5'd2};
		rom[ 1353 ] = { 5'd13,	5'd14,	5'd9,	5'd2};
		rom[ 1354 ] = { 5'd7,	5'd7,	5'd3,	5'd7};
		rom[ 1355 ] = { 5'd13,	5'd13,	5'd6,	5'd3};
		rom[ 1356 ] = { 5'd10,	5'd7,	5'd4,	5'd9};
		rom[ 1357 ] = { 5'd12,	5'd12,	5'd3,	5'd6};
		rom[ 1358 ] = { 5'd0,	5'd7,	5'd4,	5'd5};
		rom[ 1359 ] = { 5'd11,	5'd0,	5'd3,	5'd6};
		rom[ 1360 ] = { 5'd2,	5'd12,	5'd12,	5'd3};
		rom[ 1361 ] = { 5'd13,	5'd13,	5'd6,	5'd3};
		rom[ 1362 ] = { 5'd5,	5'd13,	5'd6,	5'd3};
		rom[ 1363 ] = { 5'd9,	5'd17,	5'd9,	5'd2};
		rom[ 1364 ] = { 5'd5,	5'd19,	5'd12,	5'd3};
		rom[ 1365 ] = { 5'd3,	5'd3,	5'd20,	5'd1};
		rom[ 1366 ] = { 5'd6,	5'd5,	5'd4,	5'd6};
		rom[ 1367 ] = { 5'd12,	5'd0,	5'd1,	5'd24};
		rom[ 1368 ] = { 5'd8,	5'd16,	5'd5,	5'd4};
		rom[ 1369 ] = { 5'd9,	5'd18,	5'd6,	5'd6};
		rom[ 1370 ] = { 5'd1,	5'd15,	5'd6,	5'd4};
		rom[ 1371 ] = { 5'd19,	5'd10,	5'd4,	5'd7};
		rom[ 1372 ] = { 5'd1,	5'd9,	5'd4,	5'd7};
		rom[ 1373 ] = { 5'd9,	5'd16,	5'd9,	5'd5};
		rom[ 1374 ] = { 5'd6,	5'd9,	5'd12,	5'd2};
		rom[ 1375 ] = { 5'd12,	5'd15,	5'd2,	5'd9};
		rom[ 1376 ] = { 5'd10,	5'd8,	5'd3,	5'd7};
		rom[ 1377 ] = { 5'd14,	5'd4,	5'd4,	5'd5};
		rom[ 1378 ] = { 5'd4,	5'd9,	5'd6,	5'd3};
		rom[ 1379 ] = { 5'd8,	5'd6,	5'd8,	5'd12};
		rom[ 1380 ] = { 5'd6,	5'd7,	5'd3,	5'd14};
		rom[ 1381 ] = { 5'd19,	5'd12,	5'd5,	5'd4};
		rom[ 1382 ] = { 5'd0,	5'd12,	5'd5,	5'd4};
		rom[ 1383 ] = { 5'd17,	5'd6,	5'd6,	5'd3};
		rom[ 1384 ] = { 5'd1,	5'd6,	5'd6,	5'd3};
		rom[ 1385 ] = { 5'd18,	5'd5,	5'd6,	5'd3};
		rom[ 1386 ] = { 5'd0,	5'd5,	5'd6,	5'd3};
		rom[ 1387 ] = { 5'd3,	5'd5,	5'd18,	5'd2};
		rom[ 1388 ] = { 5'd2,	5'd5,	5'd9,	5'd2};
		rom[ 1389 ] = { 5'd14,	5'd3,	5'd5,	5'd4};
		rom[ 1390 ] = { 5'd5,	5'd3,	5'd5,	5'd4};
		rom[ 1391 ] = { 5'd10,	5'd11,	5'd3,	5'd12};
		rom[ 1392 ] = { 5'd11,	5'd11,	5'd3,	5'd11};
		rom[ 1393 ] = { 5'd7,	5'd8,	5'd5,	5'd4};
		rom[ 1394 ] = { 5'd12,	5'd6,	5'd3,	5'd7};
		rom[ 1395 ] = { 5'd5,	5'd19,	5'd18,	5'd1};
		rom[ 1396 ] = { 5'd10,	5'd4,	5'd2,	5'd9};
		rom[ 1397 ] = { 5'd11,	5'd1,	5'd3,	5'd7};
		rom[ 1398 ] = { 5'd9,	5'd11,	5'd3,	5'd6};
		rom[ 1399 ] = { 5'd14,	5'd12,	5'd2,	5'd11};
		rom[ 1400 ] = { 5'd8,	5'd12,	5'd2,	5'd11};
		rom[ 1401 ] = { 5'd12,	5'd0,	5'd4,	5'd18};
		rom[ 1402 ] = { 5'd7,	5'd12,	5'd5,	5'd5};
		rom[ 1403 ] = { 5'd2,	5'd21,	5'd22,	5'd1};
		rom[ 1404 ] = { 5'd1,	5'd4,	5'd1,	5'd20};
		rom[ 1405 ] = { 5'd8,	5'd2,	5'd8,	5'd4};
		rom[ 1406 ] = { 5'd7,	5'd10,	5'd10,	5'd2};
		rom[ 1407 ] = { 5'd6,	5'd7,	5'd4,	5'd5};
		rom[ 1408 ] = { 5'd17,	5'd0,	5'd3,	5'd7};
		rom[ 1409 ] = { 5'd4,	5'd15,	5'd5,	5'd4};
		rom[ 1410 ] = { 5'd2,	5'd3,	5'd20,	5'd3};
		rom[ 1411 ] = { 5'd6,	5'd7,	5'd6,	5'd4};
		rom[ 1412 ] = { 5'd9,	5'd20,	5'd6,	5'd3};
		rom[ 1413 ] = { 5'd7,	5'd12,	5'd10,	5'd2};
		rom[ 1414 ] = { 5'd10,	5'd5,	5'd4,	5'd9};
		rom[ 1415 ] = { 5'd8,	5'd11,	5'd3,	5'd8};
		rom[ 1416 ] = { 5'd18,	5'd4,	5'd2,	5'd17};
		rom[ 1417 ] = { 5'd3,	5'd0,	5'd3,	5'd6};
		rom[ 1418 ] = { 5'd18,	5'd4,	5'd2,	5'd17};
		rom[ 1419 ] = { 5'd4,	5'd4,	5'd2,	5'd17};
		rom[ 1420 ] = { 5'd5,	5'd19,	5'd19,	5'd1};
		rom[ 1421 ] = { 5'd11,	5'd9,	5'd2,	5'd9};
		rom[ 1422 ] = { 5'd15,	5'd13,	5'd2,	5'd9};
		rom[ 1423 ] = { 5'd7,	5'd13,	5'd2,	5'd9};
		rom[ 1424 ] = { 5'd12,	5'd11,	5'd5,	5'd4};
		rom[ 1425 ] = { 5'd12,	5'd6,	5'd2,	5'd9};
		rom[ 1426 ] = { 5'd12,	5'd0,	5'd2,	5'd9};
		rom[ 1427 ] = { 5'd2,	5'd9,	5'd8,	5'd4};
		rom[ 1428 ] = { 5'd14,	5'd18,	5'd6,	5'd3};
		rom[ 1429 ] = { 5'd10,	5'd7,	5'd2,	5'd9};
		rom[ 1430 ] = { 5'd14,	5'd18,	5'd6,	5'd3};
		rom[ 1431 ] = { 5'd3,	5'd14,	5'd12,	5'd2};
		rom[ 1432 ] = { 5'd14,	5'd14,	5'd9,	5'd2};
		rom[ 1433 ] = { 5'd1,	5'd14,	5'd9,	5'd2};
		rom[ 1434 ] = { 5'd3,	5'd8,	5'd18,	5'd1};
		rom[ 1435 ] = { 5'd1,	5'd9,	5'd22,	5'd2};
		rom[ 1436 ] = { 5'd18,	5'd7,	5'd6,	5'd3};
		rom[ 1437 ] = { 5'd0,	5'd7,	5'd6,	5'd3};
		rom[ 1438 ] = { 5'd5,	5'd14,	5'd16,	5'd3};
		rom[ 1439 ] = { 5'd6,	5'd18,	5'd9,	5'd2};
		rom[ 1440 ] = { 5'd14,	5'd18,	5'd6,	5'd3};
		rom[ 1441 ] = { 5'd4,	5'd18,	5'd6,	5'd3};
		rom[ 1442 ] = { 5'd17,	5'd1,	5'd2,	5'd23};
		rom[ 1443 ] = { 5'd8,	5'd21,	5'd8,	5'd3};
		rom[ 1444 ] = { 5'd8,	5'd20,	5'd8,	5'd4};
		rom[ 1445 ] = { 5'd5,	5'd1,	5'd2,	5'd23};
		rom[ 1446 ] = { 5'd3,	5'd18,	5'd18,	5'd1};
		rom[ 1447 ] = { 5'd0,	5'd17,	5'd18,	5'd1};
		rom[ 1448 ] = { 5'd12,	5'd16,	5'd11,	5'd2};
		rom[ 1449 ] = { 5'd0,	5'd18,	5'd9,	5'd2};
		rom[ 1450 ] = { 5'd9,	5'd10,	5'd7,	5'd3};
		rom[ 1451 ] = { 5'd2,	5'd18,	5'd6,	5'd3};
		rom[ 1452 ] = { 5'd0,	5'd7,	5'd24,	5'd2};
		rom[ 1453 ] = { 5'd10,	5'd7,	5'd4,	5'd5};
		rom[ 1454 ] = { 5'd10,	5'd13,	5'd6,	5'd6};
		rom[ 1455 ] = { 5'd8,	5'd6,	5'd2,	5'd9};
		rom[ 1456 ] = { 5'd13,	5'd0,	5'd2,	5'd9};
		rom[ 1457 ] = { 5'd11,	5'd7,	5'd2,	5'd9};
		rom[ 1458 ] = { 5'd2,	5'd2,	5'd20,	5'd1};
		rom[ 1459 ] = { 5'd1,	5'd18,	5'd6,	5'd3};
		rom[ 1460 ] = { 5'd13,	5'd2,	5'd2,	5'd13};
		rom[ 1461 ] = { 5'd12,	5'd7,	5'd6,	5'd4};
		rom[ 1462 ] = { 5'd10,	5'd1,	5'd2,	5'd13};
		rom[ 1463 ] = { 5'd7,	5'd0,	5'd1,	5'd18};
		rom[ 1464 ] = { 5'd14,	5'd3,	5'd5,	5'd5};
		rom[ 1465 ] = { 5'd10,	5'd15,	5'd4,	5'd8};
		rom[ 1466 ] = { 5'd11,	5'd10,	5'd2,	5'd9};
		rom[ 1467 ] = { 5'd10,	5'd3,	5'd2,	5'd9};
		rom[ 1468 ] = { 5'd20,	5'd0,	5'd3,	5'd7};
		rom[ 1469 ] = { 5'd1,	5'd0,	5'd3,	5'd7};
		rom[ 1470 ] = { 5'd17,	5'd0,	5'd3,	5'd8};
		rom[ 1471 ] = { 5'd9,	5'd4,	5'd2,	5'd10};
		rom[ 1472 ] = { 5'd12,	5'd17,	5'd9,	5'd3};
		rom[ 1473 ] = { 5'd12,	5'd20,	5'd11,	5'd4};
		rom[ 1474 ] = { 5'd14,	5'd3,	5'd5,	5'd5};
		rom[ 1475 ] = { 5'd5,	5'd3,	5'd5,	5'd5};
		rom[ 1476 ] = { 5'd16,	5'd6,	5'd4,	5'd16};
		rom[ 1477 ] = { 5'd4,	5'd6,	5'd4,	5'd16};
		rom[ 1478 ] = { 5'd10,	5'd14,	5'd5,	5'd5};
		rom[ 1479 ] = { 5'd1,	5'd19,	5'd21,	5'd1};
		rom[ 1480 ] = { 5'd15,	5'd2,	5'd9,	5'd2};
		rom[ 1481 ] = { 5'd12,	5'd1,	5'd6,	5'd4};
		rom[ 1482 ] = { 5'd12,	5'd0,	5'd6,	5'd6};
		rom[ 1483 ] = { 5'd8,	5'd10,	5'd4,	5'd6};
		rom[ 1484 ] = { 5'd19,	5'd16,	5'd5,	5'd4};
		rom[ 1485 ] = { 5'd0,	5'd16,	5'd5,	5'd4};
		rom[ 1486 ] = { 5'd14,	5'd12,	5'd4,	5'd5};
		rom[ 1487 ] = { 5'd6,	5'd16,	5'd5,	5'd4};
		rom[ 1488 ] = { 5'd13,	5'd6,	5'd6,	5'd3};
		rom[ 1489 ] = { 5'd9,	5'd6,	5'd2,	5'd9};
		rom[ 1490 ] = { 5'd13,	5'd9,	5'd3,	5'd7};
		rom[ 1491 ] = { 5'd8,	5'd9,	5'd3,	5'd7};
		rom[ 1492 ] = { 5'd7,	5'd10,	5'd11,	5'd6};
		rom[ 1493 ] = { 5'd4,	5'd8,	5'd3,	5'd8};
		rom[ 1494 ] = { 5'd17,	5'd10,	5'd4,	5'd7};
		rom[ 1495 ] = { 5'd3,	5'd10,	5'd4,	5'd7};
		rom[ 1496 ] = { 5'd14,	5'd1,	5'd4,	5'd9};
		rom[ 1497 ] = { 5'd2,	5'd5,	5'd8,	5'd4};
		rom[ 1498 ] = { 5'd3,	5'd10,	5'd18,	5'd4};
		rom[ 1499 ] = { 5'd4,	5'd14,	5'd16,	5'd4};
		rom[ 1500 ] = { 5'd19,	5'd4,	5'd4,	5'd10};
		rom[ 1501 ] = { 5'd10,	5'd2,	5'd3,	5'd6};
		rom[ 1502 ] = { 5'd19,	5'd4,	5'd4,	5'd10};
		rom[ 1503 ] = { 5'd1,	5'd4,	5'd4,	5'd10};
		rom[ 1504 ] = { 5'd15,	5'd8,	5'd4,	5'd7};
		rom[ 1505 ] = { 5'd5,	5'd8,	5'd4,	5'd7};
		rom[ 1506 ] = { 5'd10,	5'd17,	5'd5,	5'd4};
		rom[ 1507 ] = { 5'd4,	5'd16,	5'd7,	5'd3};
		rom[ 1508 ] = { 5'd0,	5'd18,	5'd24,	5'd5};
		rom[ 1509 ] = { 5'd8,	5'd2,	5'd4,	5'd11};
		rom[ 1510 ] = { 5'd14,	5'd2,	5'd4,	5'd8};
		rom[ 1511 ] = { 5'd0,	5'd2,	5'd12,	5'd3};
		rom[ 1512 ] = { 5'd6,	5'd3,	5'd12,	5'd3};
		rom[ 1513 ] = { 5'd1,	5'd2,	5'd6,	5'd6};
		rom[ 1514 ] = { 5'd18,	5'd8,	5'd6,	5'd3};
		rom[ 1515 ] = { 5'd4,	5'd3,	5'd4,	5'd5};
		rom[ 1516 ] = { 5'd6,	5'd22,	5'd18,	5'd1};
		rom[ 1517 ] = { 5'd1,	5'd11,	5'd18,	5'd1};
		rom[ 1518 ] = { 5'd1,	5'd11,	5'd22,	5'd1};
		rom[ 1519 ] = { 5'd2,	5'd11,	5'd12,	5'd3};
		rom[ 1520 ] = { 5'd18,	5'd8,	5'd6,	5'd3};
		rom[ 1521 ] = { 5'd0,	5'd8,	5'd6,	5'd3};
		rom[ 1522 ] = { 5'd12,	5'd15,	5'd2,	5'd9};
		rom[ 1523 ] = { 5'd7,	5'd15,	5'd9,	5'd2};
		rom[ 1524 ] = { 5'd9,	5'd14,	5'd7,	5'd6};
		rom[ 1525 ] = { 5'd7,	5'd13,	5'd3,	5'd6};
		rom[ 1526 ] = { 5'd12,	5'd15,	5'd6,	5'd4};
		rom[ 1527 ] = { 5'd7,	5'd4,	5'd2,	5'd16};
		rom[ 1528 ] = { 5'd12,	5'd15,	5'd2,	5'd9};
		rom[ 1529 ] = { 5'd10,	5'd15,	5'd2,	5'd9};
		rom[ 1530 ] = { 5'd15,	5'd11,	5'd6,	5'd5};
		rom[ 1531 ] = { 5'd3,	5'd8,	5'd14,	5'd2};
		rom[ 1532 ] = { 5'd4,	5'd6,	5'd17,	5'd4};
		rom[ 1533 ] = { 5'd6,	5'd9,	5'd12,	5'd7};
		rom[ 1534 ] = { 5'd8,	5'd4,	5'd9,	5'd3};
		rom[ 1535 ] = { 5'd12,	5'd7,	5'd12,	5'd3};
		rom[ 1536 ] = { 5'd11,	5'd11,	5'd9,	5'd5};
		rom[ 1537 ] = { 5'd2,	5'd12,	5'd18,	5'd1};
		rom[ 1538 ] = { 5'd8,	5'd18,	5'd9,	5'd2};
		rom[ 1539 ] = { 5'd0,	5'd2,	5'd9,	5'd2};
		rom[ 1540 ] = { 5'd0,	5'd13,	5'd24,	5'd2};
		rom[ 1541 ] = { 5'd2,	5'd12,	5'd20,	5'd3};
		rom[ 1542 ] = { 5'd12,	5'd5,	5'd8,	5'd6};
		rom[ 1543 ] = { 5'd10,	5'd7,	5'd4,	5'd5};
		rom[ 1544 ] = { 5'd7,	5'd5,	5'd10,	5'd2};
		rom[ 1545 ] = { 5'd9,	5'd19,	5'd6,	5'd4};
		rom[ 1546 ] = { 5'd17,	5'd5,	5'd7,	5'd5};
		rom[ 1547 ] = { 5'd0,	5'd5,	5'd7,	5'd5};
		rom[ 1548 ] = { 5'd19,	5'd1,	5'd3,	5'd6};
		rom[ 1549 ] = { 5'd1,	5'd4,	5'd19,	5'd4};
		rom[ 1550 ] = { 5'd12,	5'd4,	5'd9,	5'd2};
		rom[ 1551 ] = { 5'd3,	5'd4,	5'd9,	5'd2};
		rom[ 1552 ] = { 5'd12,	5'd4,	5'd10,	5'd2};
		rom[ 1553 ] = { 5'd12,	5'd4,	5'd9,	5'd2};
		rom[ 1554 ] = { 5'd12,	5'd1,	5'd2,	5'd9};
		rom[ 1555 ] = { 5'd10,	5'd1,	5'd2,	5'd9};
		rom[ 1556 ] = { 5'd14,	5'd5,	5'd4,	5'd5};
		rom[ 1557 ] = { 5'd10,	5'd4,	5'd4,	5'd13};
		rom[ 1558 ] = { 5'd13,	5'd5,	5'd3,	5'd6};
		rom[ 1559 ] = { 5'd7,	5'd5,	5'd6,	5'd3};
		rom[ 1560 ] = { 5'd7,	5'd7,	5'd10,	5'd2};
		rom[ 1561 ] = { 5'd9,	5'd0,	5'd7,	5'd5};
		rom[ 1562 ] = { 5'd0,	5'd11,	5'd9,	5'd3};
		rom[ 1563 ] = { 5'd11,	5'd6,	5'd2,	5'd9};
		rom[ 1564 ] = { 5'd3,	5'd3,	5'd3,	5'd7};
		rom[ 1565 ] = { 5'd15,	5'd18,	5'd6,	5'd3};
		rom[ 1566 ] = { 5'd2,	5'd8,	5'd10,	5'd3};
		rom[ 1567 ] = { 5'd13,	5'd4,	5'd10,	5'd2};
		rom[ 1568 ] = { 5'd4,	5'd11,	5'd5,	5'd6};
		rom[ 1569 ] = { 5'd20,	5'd4,	5'd2,	5'd9};
		rom[ 1570 ] = { 5'd8,	5'd13,	5'd8,	5'd7};
		rom[ 1571 ] = { 5'd12,	5'd1,	5'd12,	5'd3};
		rom[ 1572 ] = { 5'd2,	5'd4,	5'd2,	5'd9};
		rom[ 1573 ] = { 5'd3,	5'd7,	5'd18,	5'd1};
		rom[ 1574 ] = { 5'd3,	5'd19,	5'd16,	5'd2};
		rom[ 1575 ] = { 5'd13,	5'd9,	5'd6,	5'd3};
		rom[ 1576 ] = { 5'd5,	5'd6,	5'd7,	5'd3};
		rom[ 1577 ] = { 5'd17,	5'd5,	5'd4,	5'd5};
		rom[ 1578 ] = { 5'd2,	5'd3,	5'd20,	5'd1};
		rom[ 1579 ] = { 5'd12,	5'd2,	5'd3,	5'd6};
		rom[ 1580 ] = { 5'd10,	5'd6,	5'd2,	5'd9};
		rom[ 1581 ] = { 5'd12,	5'd3,	5'd2,	5'd11};
		rom[ 1582 ] = { 5'd10,	5'd3,	5'd2,	5'd11};
		rom[ 1583 ] = { 5'd12,	5'd3,	5'd4,	5'd5};
		rom[ 1584 ] = { 5'd12,	5'd1,	5'd1,	5'd18};
		rom[ 1585 ] = { 5'd12,	5'd2,	5'd3,	5'd6};
		rom[ 1586 ] = { 5'd0,	5'd3,	5'd19,	5'd1};
		rom[ 1587 ] = { 5'd9,	5'd16,	5'd9,	5'd2};
		rom[ 1588 ] = { 5'd7,	5'd8,	5'd6,	5'd5};
		rom[ 1589 ] = { 5'd14,	5'd0,	5'd2,	5'd9};
		rom[ 1590 ] = { 5'd8,	5'd0,	5'd2,	5'd9};
		rom[ 1591 ] = { 5'd13,	5'd11,	5'd4,	5'd5};
		rom[ 1592 ] = { 5'd1,	5'd6,	5'd18,	5'd1};
		rom[ 1593 ] = { 5'd9,	5'd9,	5'd14,	5'd2};
		rom[ 1594 ] = { 5'd2,	5'd17,	5'd18,	5'd1};
		rom[ 1595 ] = { 5'd15,	5'd19,	5'd9,	5'd2};
		rom[ 1596 ] = { 5'd0,	5'd8,	5'd6,	5'd3};
		rom[ 1597 ] = { 5'd9,	5'd17,	5'd7,	5'd4};
		rom[ 1598 ] = { 5'd2,	5'd18,	5'd20,	5'd1};
		rom[ 1599 ] = { 5'd15,	5'd19,	5'd9,	5'd2};
		rom[ 1600 ] = { 5'd4,	5'd2,	5'd15,	5'd2};
		rom[ 1601 ] = { 5'd17,	5'd5,	5'd6,	5'd3};
		rom[ 1602 ] = { 5'd0,	5'd6,	5'd6,	5'd3};
		rom[ 1603 ] = { 5'd15,	5'd19,	5'd9,	5'd2};
		rom[ 1604 ] = { 5'd0,	5'd19,	5'd9,	5'd2};
		rom[ 1605 ] = { 5'd15,	5'd18,	5'd6,	5'd3};
		rom[ 1606 ] = { 5'd3,	5'd18,	5'd6,	5'd3};
		rom[ 1607 ] = { 5'd20,	5'd13,	5'd4,	5'd5};
		rom[ 1608 ] = { 5'd8,	5'd14,	5'd8,	5'd4};
		rom[ 1609 ] = { 5'd13,	5'd18,	5'd3,	5'd6};
		rom[ 1610 ] = { 5'd0,	5'd13,	5'd4,	5'd5};
		rom[ 1611 ] = { 5'd0,	5'd17,	5'd24,	5'd3};
		rom[ 1612 ] = { 5'd5,	5'd2,	5'd6,	5'd4};
		rom[ 1613 ] = { 5'd11,	5'd9,	5'd3,	5'd6};
		rom[ 1614 ] = { 5'd4,	5'd5,	5'd16,	5'd2};
		rom[ 1615 ] = { 5'd10,	5'd7,	5'd4,	5'd5};
		rom[ 1616 ] = { 5'd8,	5'd8,	5'd5,	5'd4};
		rom[ 1617 ] = { 5'd11,	5'd9,	5'd9,	5'd4};
		rom[ 1618 ] = { 5'd4,	5'd9,	5'd9,	5'd4};
		rom[ 1619 ] = { 5'd14,	5'd9,	5'd6,	5'd3};
		rom[ 1620 ] = { 5'd2,	5'd8,	5'd20,	5'd4};
		rom[ 1621 ] = { 5'd4,	5'd12,	5'd17,	5'd8};
		rom[ 1622 ] = { 5'd8,	5'd10,	5'd7,	5'd3};
		rom[ 1623 ] = { 5'd1,	5'd10,	5'd23,	5'd1};
		rom[ 1624 ] = { 5'd9,	5'd0,	5'd2,	5'd9};
		rom[ 1625 ] = { 5'd13,	5'd3,	5'd2,	5'd9};
		rom[ 1626 ] = { 5'd10,	5'd1,	5'd2,	5'd13};
		rom[ 1627 ] = { 5'd4,	5'd23,	5'd18,	5'd1};
		rom[ 1628 ] = { 5'd6,	5'd10,	5'd3,	5'd6};
		rom[ 1629 ] = { 5'd14,	5'd0,	5'd1,	5'd24};
		rom[ 1630 ] = { 5'd9,	5'd0,	5'd1,	5'd24};
		rom[ 1631 ] = { 5'd9,	5'd2,	5'd6,	5'd10};
		rom[ 1632 ] = { 5'd9,	5'd13,	5'd5,	5'd6};
		rom[ 1633 ] = { 5'd9,	5'd21,	5'd6,	5'd3};
		rom[ 1634 ] = { 5'd11,	5'd1,	5'd2,	5'd11};
		rom[ 1635 ] = { 5'd9,	5'd7,	5'd5,	5'd4};
		rom[ 1636 ] = { 5'd12,	5'd0,	5'd5,	5'd18};
		rom[ 1637 ] = { 5'd14,	5'd1,	5'd2,	5'd16};
		rom[ 1638 ] = { 5'd8,	5'd1,	5'd2,	5'd16};
		rom[ 1639 ] = { 5'd18,	5'd5,	5'd6,	5'd3};
		rom[ 1640 ] = { 5'd3,	5'd6,	5'd18,	5'd1};
		rom[ 1641 ] = { 5'd18,	5'd5,	5'd6,	5'd3};
		rom[ 1642 ] = { 5'd0,	5'd5,	5'd6,	5'd3};
		rom[ 1643 ] = { 5'd13,	5'd13,	5'd11,	5'd2};
		rom[ 1644 ] = { 5'd10,	5'd7,	5'd5,	5'd4};
		rom[ 1645 ] = { 5'd11,	5'd9,	5'd5,	5'd7};
		rom[ 1646 ] = { 5'd8,	5'd9,	5'd5,	5'd7};
		rom[ 1647 ] = { 5'd16,	5'd4,	5'd3,	5'd6};
		rom[ 1648 ] = { 5'd5,	5'd6,	5'd5,	5'd4};
		rom[ 1649 ] = { 5'd7,	5'd21,	5'd8,	5'd3};
		rom[ 1650 ] = { 5'd9,	5'd21,	5'd8,	5'd3};
		rom[ 1651 ] = { 5'd13,	5'd5,	5'd11,	5'd7};
		rom[ 1652 ] = { 5'd3,	5'd10,	5'd4,	5'd5};
		rom[ 1653 ] = { 5'd20,	5'd0,	5'd3,	5'd6};
		rom[ 1654 ] = { 5'd7,	5'd2,	5'd2,	5'd18};
		rom[ 1655 ] = { 5'd15,	5'd0,	5'd2,	5'd9};
		rom[ 1656 ] = { 5'd0,	5'd15,	5'd7,	5'd3};
		rom[ 1657 ] = { 5'd19,	5'd13,	5'd4,	5'd5};
		rom[ 1658 ] = { 5'd1,	5'd0,	5'd3,	5'd6};
		rom[ 1659 ] = { 5'd12,	5'd7,	5'd3,	5'd6};
		rom[ 1660 ] = { 5'd1,	5'd13,	5'd4,	5'd5};
		rom[ 1661 ] = { 5'd3,	5'd22,	5'd19,	5'd1};
		rom[ 1662 ] = { 5'd8,	5'd3,	5'd2,	5'd13};
		rom[ 1663 ] = { 5'd5,	5'd11,	5'd18,	5'd1};
		rom[ 1664 ] = { 5'd9,	5'd7,	5'd5,	5'd4};
		rom[ 1665 ] = { 5'd11,	5'd7,	5'd4,	5'd5};
		rom[ 1666 ] = { 5'd4,	5'd3,	5'd16,	5'd2};
		rom[ 1667 ] = { 5'd6,	5'd1,	5'd18,	5'd1};
		rom[ 1668 ] = { 5'd5,	5'd1,	5'd5,	5'd4};
		rom[ 1669 ] = { 5'd17,	5'd18,	5'd6,	5'd3};
		rom[ 1670 ] = { 5'd11,	5'd15,	5'd6,	5'd3};
		rom[ 1671 ] = { 5'd1,	5'd10,	5'd11,	5'd4};
		rom[ 1672 ] = { 5'd10,	5'd9,	5'd3,	5'd6};
		rom[ 1673 ] = { 5'd10,	5'd11,	5'd4,	5'd5};
		rom[ 1674 ] = { 5'd11,	5'd7,	5'd5,	5'd7};
		rom[ 1675 ] = { 5'd11,	5'd2,	5'd4,	5'd10};
		rom[ 1676 ] = { 5'd9,	5'd2,	5'd4,	5'd10};
		rom[ 1677 ] = { 5'd15,	5'd4,	5'd9,	5'd3};
		rom[ 1678 ] = { 5'd0,	5'd8,	5'd10,	5'd3};
		rom[ 1679 ] = { 5'd2,	5'd9,	5'd21,	5'd2};
		rom[ 1680 ] = { 5'd0,	5'd4,	5'd11,	5'd8};
		rom[ 1681 ] = { 5'd9,	5'd11,	5'd6,	5'd11};
		rom[ 1682 ] = { 5'd9,	5'd7,	5'd3,	5'd6};
		rom[ 1683 ] = { 5'd18,	5'd0,	5'd6,	5'd9};
		rom[ 1684 ] = { 5'd0,	5'd0,	5'd6,	5'd9};
		rom[ 1685 ] = { 5'd12,	5'd1,	5'd11,	5'd2};
		rom[ 1686 ] = { 5'd3,	5'd2,	5'd18,	5'd2};
		rom[ 1687 ] = { 5'd2,	5'd7,	5'd22,	5'd2};
		rom[ 1688 ] = { 5'd5,	5'd3,	5'd6,	5'd3};
		rom[ 1689 ] = { 5'd12,	5'd14,	5'd2,	5'd9};
		rom[ 1690 ] = { 5'd10,	5'd14,	5'd2,	5'd9};
		rom[ 1691 ] = { 5'd5,	5'd19,	5'd18,	5'd1};
		rom[ 1692 ] = { 5'd9,	5'd0,	5'd3,	5'd13};
		rom[ 1693 ] = { 5'd7,	5'd4,	5'd6,	5'd4};
		rom[ 1694 ] = { 5'd9,	5'd2,	5'd4,	5'd6};
		rom[ 1695 ] = { 5'd4,	5'd2,	5'd18,	5'd1};
		rom[ 1696 ] = { 5'd0,	5'd12,	5'd6,	5'd4};
		rom[ 1697 ] = { 5'd11,	5'd15,	5'd2,	5'd9};
		rom[ 1698 ] = { 5'd11,	5'd10,	5'd2,	5'd13};
		rom[ 1699 ] = { 5'd6,	5'd18,	5'd18,	5'd1};
		rom[ 1700 ] = { 5'd11,	5'd4,	5'd2,	5'd9};
		rom[ 1701 ] = { 5'd12,	5'd0,	5'd2,	5'd9};
		rom[ 1702 ] = { 5'd5,	5'd6,	5'd5,	5'd4};
		rom[ 1703 ] = { 5'd14,	5'd13,	5'd5,	5'd4};
		rom[ 1704 ] = { 5'd5,	5'd13,	5'd5,	5'd4};
		rom[ 1705 ] = { 5'd14,	5'd13,	5'd9,	5'd2};
		rom[ 1706 ] = { 5'd0,	5'd7,	5'd23,	5'd5};
		rom[ 1707 ] = { 5'd16,	5'd6,	5'd8,	5'd6};
		rom[ 1708 ] = { 5'd4,	5'd18,	5'd6,	5'd3};
		rom[ 1709 ] = { 5'd8,	5'd20,	5'd9,	5'd2};
		rom[ 1710 ] = { 5'd0,	5'd18,	5'd18,	5'd1};
		rom[ 1711 ] = { 5'd13,	5'd13,	5'd11,	5'd2};
		rom[ 1712 ] = { 5'd0,	5'd13,	5'd11,	5'd2};
		rom[ 1713 ] = { 5'd12,	5'd9,	5'd12,	5'd3};
		rom[ 1714 ] = { 5'd6,	5'd20,	5'd8,	5'd4};
		rom[ 1715 ] = { 5'd10,	5'd18,	5'd14,	5'd2};
		rom[ 1716 ] = { 5'd1,	5'd2,	5'd21,	5'd1};
		rom[ 1717 ] = { 5'd0,	5'd2,	5'd12,	5'd3};
		rom[ 1718 ] = { 5'd6,	5'd15,	5'd4,	5'd5};
		rom[ 1719 ] = { 5'd9,	5'd11,	5'd7,	5'd3};
		rom[ 1720 ] = { 5'd1,	5'd18,	5'd6,	5'd3};
		rom[ 1721 ] = { 5'd10,	5'd19,	5'd4,	5'd5};
		rom[ 1722 ] = { 5'd7,	5'd12,	5'd4,	5'd5};
		rom[ 1723 ] = { 5'd9,	5'd12,	5'd6,	5'd4};
		rom[ 1724 ] = { 5'd10,	5'd1,	5'd3,	5'd6};
		rom[ 1725 ] = { 5'd3,	5'd15,	5'd19,	5'd1};
		rom[ 1726 ] = { 5'd7,	5'd7,	5'd5,	5'd5};
		rom[ 1727 ] = { 5'd3,	5'd12,	5'd9,	5'd12};
		rom[ 1728 ] = { 5'd10,	5'd0,	5'd2,	5'd12};
		rom[ 1729 ] = { 5'd3,	5'd3,	5'd17,	5'd3};
		rom[ 1730 ] = { 5'd10,	5'd0,	5'd4,	5'd11};
		rom[ 1731 ] = { 5'd4,	5'd0,	5'd3,	5'd13};
		rom[ 1732 ] = { 5'd5,	5'd11,	5'd16,	5'd3};
		rom[ 1733 ] = { 5'd8,	5'd14,	5'd5,	5'd6};
		rom[ 1734 ] = { 5'd9,	5'd21,	5'd6,	5'd3};
		rom[ 1735 ] = { 5'd3,	5'd0,	5'd3,	5'd6};
		rom[ 1736 ] = { 5'd2,	5'd1,	5'd20,	5'd1};
		rom[ 1737 ] = { 5'd9,	5'd6,	5'd5,	5'd10};
		rom[ 1738 ] = { 5'd11,	5'd6,	5'd2,	5'd9};
		rom[ 1739 ] = { 5'd11,	5'd0,	5'd2,	5'd9};
		rom[ 1740 ] = { 5'd16,	5'd0,	5'd2,	5'd9};
		rom[ 1741 ] = { 5'd7,	5'd18,	5'd9,	5'd2};
		rom[ 1742 ] = { 5'd16,	5'd0,	5'd2,	5'd9};
		rom[ 1743 ] = { 5'd6,	5'd0,	5'd2,	5'd9};
		rom[ 1744 ] = { 5'd19,	5'd1,	5'd2,	5'd16};
		rom[ 1745 ] = { 5'd3,	5'd1,	5'd2,	5'd16};
		rom[ 1746 ] = { 5'd14,	5'd16,	5'd6,	5'd3};
		rom[ 1747 ] = { 5'd0,	5'd3,	5'd6,	5'd3};
		rom[ 1748 ] = { 5'd9,	5'd5,	5'd3,	5'd6};
		rom[ 1749 ] = { 5'd6,	5'd10,	5'd3,	5'd6};
		rom[ 1750 ] = { 5'd14,	5'd15,	5'd3,	5'd8};
		rom[ 1751 ] = { 5'd4,	5'd10,	5'd7,	5'd6};
		rom[ 1752 ] = { 5'd7,	5'd8,	5'd12,	5'd2};
		rom[ 1753 ] = { 5'd9,	5'd2,	5'd2,	5'd20};
		rom[ 1754 ] = { 5'd14,	5'd16,	5'd6,	5'd3};
		rom[ 1755 ] = { 5'd12,	5'd6,	5'd2,	5'd9};
		rom[ 1756 ] = { 5'd14,	5'd16,	5'd6,	5'd3};
		rom[ 1757 ] = { 5'd5,	5'd22,	5'd14,	5'd2};
		rom[ 1758 ] = { 5'd4,	5'd10,	5'd16,	5'd6};
		rom[ 1759 ] = { 5'd11,	5'd6,	5'd2,	5'd9};
		rom[ 1760 ] = { 5'd3,	5'd2,	5'd21,	5'd2};
		rom[ 1761 ] = { 5'd4,	5'd16,	5'd6,	5'd3};
		rom[ 1762 ] = { 5'd16,	5'd20,	5'd5,	5'd4};
		rom[ 1763 ] = { 5'd4,	5'd0,	5'd8,	5'd8};
		rom[ 1764 ] = { 5'd13,	5'd6,	5'd7,	5'd3};
		rom[ 1765 ] = { 5'd10,	5'd10,	5'd4,	5'd5};
		rom[ 1766 ] = { 5'd15,	5'd15,	5'd6,	5'd4};
		rom[ 1767 ] = { 5'd12,	5'd7,	5'd6,	5'd4};
		rom[ 1768 ] = { 5'd12,	5'd6,	5'd7,	5'd3};
		rom[ 1769 ] = { 5'd3,	5'd6,	5'd9,	5'd5};
		rom[ 1770 ] = { 5'd12,	5'd0,	5'd6,	5'd21};
		rom[ 1771 ] = { 5'd8,	5'd0,	5'd8,	5'd21};
		rom[ 1772 ] = { 5'd6,	5'd19,	5'd18,	5'd1};
		rom[ 1773 ] = { 5'd0,	5'd17,	5'd9,	5'd2};
		rom[ 1774 ] = { 5'd4,	5'd4,	5'd19,	5'd1};
		rom[ 1775 ] = { 5'd0,	5'd4,	5'd24,	5'd1};
		rom[ 1776 ] = { 5'd15,	5'd16,	5'd9,	5'd2};
		rom[ 1777 ] = { 5'd0,	5'd16,	5'd9,	5'd2};
		rom[ 1778 ] = { 5'd6,	5'd16,	5'd18,	5'd1};
		rom[ 1779 ] = { 5'd3,	5'd18,	5'd18,	5'd1};
		rom[ 1780 ] = { 5'd13,	5'd0,	5'd1,	5'd23};
		rom[ 1781 ] = { 5'd6,	5'd3,	5'd8,	5'd3};
		rom[ 1782 ] = { 5'd6,	5'd17,	5'd18,	5'd1};
		rom[ 1783 ] = { 5'd10,	5'd0,	5'd1,	5'd23};
		rom[ 1784 ] = { 5'd10,	5'd12,	5'd4,	5'd5};
		rom[ 1785 ] = { 5'd7,	5'd12,	5'd10,	5'd4};
		rom[ 1786 ] = { 5'd17,	5'd9,	5'd3,	5'd7};
		rom[ 1787 ] = { 5'd2,	5'd3,	5'd10,	5'd3};
		rom[ 1788 ] = { 5'd11,	5'd7,	5'd5,	5'd6};
		rom[ 1789 ] = { 5'd1,	5'd4,	5'd6,	5'd5};
		rom[ 1790 ] = { 5'd15,	5'd3,	5'd9,	5'd2};
		rom[ 1791 ] = { 5'd1,	5'd2,	5'd4,	5'd5};
		rom[ 1792 ] = { 5'd10,	5'd5,	5'd5,	5'd4};
		rom[ 1793 ] = { 5'd11,	5'd0,	5'd7,	5'd24};
		rom[ 1794 ] = { 5'd7,	5'd19,	5'd10,	5'd2};
		rom[ 1795 ] = { 5'd10,	5'd19,	5'd4,	5'd5};
		rom[ 1796 ] = { 5'd15,	5'd15,	5'd2,	5'd9};
		rom[ 1797 ] = { 5'd3,	5'd22,	5'd18,	5'd1};
		rom[ 1798 ] = { 5'd15,	5'd15,	5'd2,	5'd9};
		rom[ 1799 ] = { 5'd7,	5'd15,	5'd2,	5'd9};
		rom[ 1800 ] = { 5'd12,	5'd6,	5'd2,	5'd9};
		rom[ 1801 ] = { 5'd9,	5'd3,	5'd2,	5'd11};
		rom[ 1802 ] = { 5'd15,	5'd3,	5'd9,	5'd2};
		rom[ 1803 ] = { 5'd5,	5'd8,	5'd14,	5'd4};
		rom[ 1804 ] = { 5'd8,	5'd4,	5'd15,	5'd3};
		rom[ 1805 ] = { 5'd7,	5'd2,	5'd4,	5'd5};
		rom[ 1806 ] = { 5'd12,	5'd2,	5'd3,	5'd12};
		rom[ 1807 ] = { 5'd9,	5'd2,	5'd3,	5'd12};
		rom[ 1808 ] = { 5'd7,	5'd7,	5'd6,	5'd4};
		rom[ 1809 ] = { 5'd10,	5'd3,	5'd4,	5'd10};
		rom[ 1810 ] = { 5'd13,	5'd6,	5'd8,	5'd3};
		rom[ 1811 ] = { 5'd9,	5'd1,	5'd6,	5'd9};
		rom[ 1812 ] = { 5'd9,	5'd8,	5'd6,	5'd5};
		rom[ 1813 ] = { 5'd0,	5'd0,	5'd12,	5'd11};
		rom[ 1814 ] = { 5'd14,	5'd18,	5'd9,	5'd2};
		rom[ 1815 ] = { 5'd0,	5'd20,	5'd24,	5'd4};
		rom[ 1816 ] = { 5'd12,	5'd19,	5'd11,	5'd2};
		rom[ 1817 ] = { 5'd1,	5'd18,	5'd9,	5'd2};
		rom[ 1818 ] = { 5'd7,	5'd8,	5'd5,	5'd4};
		rom[ 1819 ] = { 5'd11,	5'd15,	5'd2,	5'd9};
		rom[ 1820 ] = { 5'd16,	5'd18,	5'd6,	5'd3};
		rom[ 1821 ] = { 5'd2,	5'd18,	5'd6,	5'd3};
		rom[ 1822 ] = { 5'd8,	5'd6,	5'd16,	5'd3};
		rom[ 1823 ] = { 5'd0,	5'd7,	5'd10,	5'd2};
		rom[ 1824 ] = { 5'd5,	5'd6,	5'd18,	5'd1};
		rom[ 1825 ] = { 5'd2,	5'd9,	5'd9,	5'd3};
		rom[ 1826 ] = { 5'd14,	5'd5,	5'd10,	5'd3};
		rom[ 1827 ] = { 5'd3,	5'd7,	5'd18,	5'd1};
		rom[ 1828 ] = { 5'd9,	5'd4,	5'd15,	5'd2};
		rom[ 1829 ] = { 5'd4,	5'd10,	5'd15,	5'd2};
		rom[ 1830 ] = { 5'd12,	5'd5,	5'd12,	5'd2};
		rom[ 1831 ] = { 5'd9,	5'd8,	5'd2,	5'd12};
		rom[ 1832 ] = { 5'd13,	5'd0,	5'd2,	5'd9};
		rom[ 1833 ] = { 5'd0,	5'd12,	5'd3,	5'd6};
		rom[ 1834 ] = { 5'd14,	5'd14,	5'd10,	5'd2};
		rom[ 1835 ] = { 5'd2,	5'd10,	5'd18,	5'd3};
		rom[ 1836 ] = { 5'd11,	5'd17,	5'd10,	5'd3};
		rom[ 1837 ] = { 5'd7,	5'd6,	5'd5,	5'd4};
		rom[ 1838 ] = { 5'd13,	5'd6,	5'd7,	5'd3};
		rom[ 1839 ] = { 5'd7,	5'd13,	5'd3,	5'd7};
		rom[ 1840 ] = { 5'd17,	5'd10,	5'd3,	5'd6};
		rom[ 1841 ] = { 5'd4,	5'd10,	5'd3,	5'd6};
		rom[ 1842 ] = { 5'd13,	5'd9,	5'd4,	5'd6};
		rom[ 1843 ] = { 5'd10,	5'd3,	5'd2,	5'd14};
		rom[ 1844 ] = { 5'd18,	5'd0,	5'd1,	5'd18};
		rom[ 1845 ] = { 5'd12,	5'd12,	5'd8,	5'd12};
		rom[ 1846 ] = { 5'd17,	5'd0,	5'd2,	5'd14};
		rom[ 1847 ] = { 5'd5,	5'd0,	5'd2,	5'd14};
		rom[ 1848 ] = { 5'd16,	5'd2,	5'd4,	5'd20};
		rom[ 1849 ] = { 5'd4,	5'd2,	5'd4,	5'd20};
		rom[ 1850 ] = { 5'd18,	5'd0,	5'd2,	5'd17};
		rom[ 1851 ] = { 5'd4,	5'd0,	5'd2,	5'd17};
		rom[ 1852 ] = { 5'd15,	5'd8,	5'd9,	5'd2};
		rom[ 1853 ] = { 5'd0,	5'd8,	5'd9,	5'd2};
		rom[ 1854 ] = { 5'd20,	5'd1,	5'd2,	5'd13};
		rom[ 1855 ] = { 5'd2,	5'd1,	5'd2,	5'd13};
		rom[ 1856 ] = { 5'd16,	5'd0,	5'd2,	5'd9};
		rom[ 1857 ] = { 5'd9,	5'd10,	5'd4,	5'd7};
		rom[ 1858 ] = { 5'd12,	5'd11,	5'd12,	5'd2};
		rom[ 1859 ] = { 5'd0,	5'd11,	5'd12,	5'd2};
		rom[ 1860 ] = { 5'd5,	5'd10,	5'd14,	5'd3};
		rom[ 1861 ] = { 5'd0,	5'd16,	5'd20,	5'd1};
		rom[ 1862 ] = { 5'd12,	5'd10,	5'd4,	5'd5};
		rom[ 1863 ] = { 5'd5,	5'd7,	5'd13,	5'd3};
		rom[ 1864 ] = { 5'd10,	5'd8,	5'd6,	5'd6};
		rom[ 1865 ] = { 5'd8,	5'd0,	5'd2,	5'd9};
		rom[ 1866 ] = { 5'd6,	5'd11,	5'd12,	5'd2};
		rom[ 1867 ] = { 5'd3,	5'd6,	5'd15,	5'd4};
		rom[ 1868 ] = { 5'd16,	5'd0,	5'd4,	5'd5};
		rom[ 1869 ] = { 5'd6,	5'd15,	5'd6,	5'd3};
		rom[ 1870 ] = { 5'd8,	5'd14,	5'd8,	5'd5};
		rom[ 1871 ] = { 5'd6,	5'd1,	5'd1,	5'd18};
		rom[ 1872 ] = { 5'd10,	5'd0,	5'd2,	5'd14};
		rom[ 1873 ] = { 5'd11,	5'd3,	5'd2,	5'd9};
		rom[ 1874 ] = { 5'd14,	5'd2,	5'd6,	5'd3};
		rom[ 1875 ] = { 5'd0,	5'd6,	5'd17,	5'd2};
		rom[ 1876 ] = { 5'd16,	5'd20,	5'd5,	5'd4};
		rom[ 1877 ] = { 5'd3,	5'd20,	5'd5,	5'd4};
		rom[ 1878 ] = { 5'd6,	5'd19,	5'd18,	5'd1};
		rom[ 1879 ] = { 5'd4,	5'd0,	5'd4,	5'd5};
		rom[ 1880 ] = { 5'd17,	5'd3,	5'd3,	5'd6};
		rom[ 1881 ] = { 5'd2,	5'd12,	5'd2,	5'd12};
		rom[ 1882 ] = { 5'd2,	5'd4,	5'd21,	5'd1};
		rom[ 1883 ] = { 5'd4,	5'd3,	5'd3,	5'd6};
		rom[ 1884 ] = { 5'd18,	5'd8,	5'd6,	5'd3};
		rom[ 1885 ] = { 5'd8,	5'd15,	5'd8,	5'd9};
		rom[ 1886 ] = { 5'd6,	5'd13,	5'd9,	5'd5};
		rom[ 1887 ] = { 5'd6,	5'd6,	5'd5,	5'd6};
		rom[ 1888 ] = { 5'd14,	5'd9,	5'd3,	5'd6};
		rom[ 1889 ] = { 5'd8,	5'd0,	5'd5,	5'd11};
		rom[ 1890 ] = { 5'd15,	5'd9,	5'd3,	5'd6};
		rom[ 1891 ] = { 5'd6,	5'd9,	5'd3,	5'd6};
		rom[ 1892 ] = { 5'd14,	5'd5,	5'd5,	5'd4};
		rom[ 1893 ] = { 5'd4,	5'd4,	5'd8,	5'd4};
		rom[ 1894 ] = { 5'd7,	5'd7,	5'd6,	5'd3};
		rom[ 1895 ] = { 5'd8,	5'd0,	5'd3,	5'd13};
		rom[ 1896 ] = { 5'd13,	5'd0,	5'd2,	5'd9};
		rom[ 1897 ] = { 5'd9,	5'd0,	5'd2,	5'd9};
		rom[ 1898 ] = { 5'd8,	5'd4,	5'd10,	5'd3};
		rom[ 1899 ] = { 5'd0,	5'd3,	5'd18,	5'd1};
		rom[ 1900 ] = { 5'd17,	5'd13,	5'd7,	5'd3};
		rom[ 1901 ] = { 5'd0,	5'd13,	5'd7,	5'd3};
		rom[ 1902 ] = { 5'd21,	5'd2,	5'd1,	5'd21};
		rom[ 1903 ] = { 5'd0,	5'd13,	5'd5,	5'd4};
		rom[ 1904 ] = { 5'd12,	5'd8,	5'd12,	5'd2};
		rom[ 1905 ] = { 5'd1,	5'd9,	5'd20,	5'd1};
		rom[ 1906 ] = { 5'd5,	5'd8,	5'd19,	5'd1};
		rom[ 1907 ] = { 5'd1,	5'd14,	5'd9,	5'd2};
		rom[ 1908 ] = { 5'd6,	5'd14,	5'd14,	5'd4};
		rom[ 1909 ] = { 5'd5,	5'd12,	5'd14,	5'd6};
		rom[ 1910 ] = { 5'd14,	5'd12,	5'd3,	5'd7};
		rom[ 1911 ] = { 5'd1,	5'd17,	5'd18,	5'd2};
		rom[ 1912 ] = { 5'd11,	5'd17,	5'd6,	5'd3};
		rom[ 1913 ] = { 5'd0,	5'd8,	5'd9,	5'd2};
		rom[ 1914 ] = { 5'd13,	5'd10,	5'd10,	5'd3};
		rom[ 1915 ] = { 5'd1,	5'd10,	5'd10,	5'd3};
		rom[ 1916 ] = { 5'd0,	5'd9,	5'd12,	5'd2};
		rom[ 1917 ] = { 5'd1,	5'd12,	5'd10,	5'd4};
		rom[ 1918 ] = { 5'd14,	5'd12,	5'd3,	5'd7};
		rom[ 1919 ] = { 5'd7,	5'd12,	5'd3,	5'd7};
		rom[ 1920 ] = { 5'd12,	5'd12,	5'd4,	5'd5};
		rom[ 1921 ] = { 5'd8,	5'd12,	5'd4,	5'd5};
		rom[ 1922 ] = { 5'd13,	5'd10,	5'd2,	5'd10};
		rom[ 1923 ] = { 5'd11,	5'd15,	5'd10,	5'd2};
		rom[ 1924 ] = { 5'd9,	5'd10,	5'd3,	5'd6};
		rom[ 1925 ] = { 5'd7,	5'd1,	5'd7,	5'd3};
		rom[ 1926 ] = { 5'd6,	5'd7,	5'd13,	5'd3};
		rom[ 1927 ] = { 5'd10,	5'd5,	5'd4,	5'd5};
		rom[ 1928 ] = { 5'd10,	5'd12,	5'd10,	5'd2};
		rom[ 1929 ] = { 5'd6,	5'd16,	5'd5,	5'd4};
		rom[ 1930 ] = { 5'd15,	5'd0,	5'd2,	5'd9};
		rom[ 1931 ] = { 5'd8,	5'd10,	5'd6,	5'd6};
		rom[ 1932 ] = { 5'd11,	5'd4,	5'd9,	5'd2};
		rom[ 1933 ] = { 5'd8,	5'd20,	5'd7,	5'd3};
		rom[ 1934 ] = { 5'd1,	5'd11,	5'd22,	5'd1};
		rom[ 1935 ] = { 5'd0,	5'd18,	5'd18,	5'd1};
		rom[ 1936 ] = { 5'd15,	5'd0,	5'd2,	5'd9};
		rom[ 1937 ] = { 5'd7,	5'd0,	5'd2,	5'd9};
		rom[ 1938 ] = { 5'd20,	5'd2,	5'd2,	5'd20};
		rom[ 1939 ] = { 5'd2,	5'd2,	5'd2,	5'd20};
		rom[ 1940 ] = { 5'd14,	5'd7,	5'd3,	5'd7};
		rom[ 1941 ] = { 5'd2,	5'd1,	5'd2,	5'd9};
		rom[ 1942 ] = { 5'd12,	5'd16,	5'd9,	5'd2};
		rom[ 1943 ] = { 5'd1,	5'd15,	5'd9,	5'd2};
		rom[ 1944 ] = { 5'd7,	5'd8,	5'd15,	5'd2};
		rom[ 1945 ] = { 5'd8,	5'd8,	5'd3,	5'd6};
		rom[ 1946 ] = { 5'd12,	5'd6,	5'd6,	5'd3};
		rom[ 1947 ] = { 5'd2,	5'd19,	5'd10,	5'd2};
		rom[ 1948 ] = { 5'd14,	5'd18,	5'd6,	5'd3};
		rom[ 1949 ] = { 5'd3,	5'd5,	5'd9,	5'd7};
		rom[ 1950 ] = { 5'd17,	5'd6,	5'd2,	5'd9};
		rom[ 1951 ] = { 5'd5,	5'd6,	5'd2,	5'd9};
		rom[ 1952 ] = { 5'd13,	5'd0,	5'd2,	5'd9};
		rom[ 1953 ] = { 5'd9,	5'd0,	5'd2,	5'd9};
		rom[ 1954 ] = { 5'd13,	5'd5,	5'd2,	5'd9};
		rom[ 1955 ] = { 5'd12,	5'd5,	5'd3,	5'd6};
		rom[ 1956 ] = { 5'd12,	5'd1,	5'd8,	5'd3};
		rom[ 1957 ] = { 5'd11,	5'd13,	5'd2,	5'd11};
		rom[ 1958 ] = { 5'd20,	5'd1,	5'd3,	5'd6};
		rom[ 1959 ] = { 5'd1,	5'd18,	5'd18,	5'd1};
		rom[ 1960 ] = { 5'd7,	5'd17,	5'd10,	5'd4};
		rom[ 1961 ] = { 5'd6,	5'd20,	5'd10,	5'd2};
		rom[ 1962 ] = { 5'd9,	5'd16,	5'd9,	5'd2};
		rom[ 1963 ] = { 5'd1,	5'd1,	5'd3,	5'd6};
		rom[ 1964 ] = { 5'd19,	5'd8,	5'd5,	5'd4};
		rom[ 1965 ] = { 5'd4,	5'd0,	5'd4,	5'd8};
		rom[ 1966 ] = { 5'd3,	5'd6,	5'd19,	5'd1};
		rom[ 1967 ] = { 5'd1,	5'd5,	5'd6,	5'd3};
		rom[ 1968 ] = { 5'd9,	5'd1,	5'd7,	5'd8};
		rom[ 1969 ] = { 5'd4,	5'd5,	5'd16,	5'd4};
		rom[ 1970 ] = { 5'd6,	5'd1,	5'd18,	5'd1};
		rom[ 1971 ] = { 5'd4,	5'd11,	5'd10,	5'd7};
		rom[ 1972 ] = { 5'd15,	5'd11,	5'd4,	5'd5};
		rom[ 1973 ] = { 5'd9,	5'd18,	5'd6,	5'd3};
		rom[ 1974 ] = { 5'd12,	5'd18,	5'd4,	5'd6};
		rom[ 1975 ] = { 5'd6,	5'd15,	5'd3,	5'd9};
		rom[ 1976 ] = { 5'd15,	5'd11,	5'd6,	5'd4};
		rom[ 1977 ] = { 5'd3,	5'd11,	5'd6,	5'd4};
		rom[ 1978 ] = { 5'd14,	5'd9,	5'd9,	5'd3};
		rom[ 1979 ] = { 5'd1,	5'd15,	5'd12,	5'd2};
		rom[ 1980 ] = { 5'd14,	5'd17,	5'd10,	5'd2};
		rom[ 1981 ] = { 5'd0,	5'd17,	5'd10,	5'd2};
		rom[ 1982 ] = { 5'd15,	5'd16,	5'd6,	5'd3};
		rom[ 1983 ] = { 5'd3,	5'd16,	5'd6,	5'd3};
		rom[ 1984 ] = { 5'd9,	5'd5,	5'd4,	5'd8};
		rom[ 1985 ] = { 5'd1,	5'd18,	5'd6,	5'd3};
		rom[ 1986 ] = { 5'd13,	5'd21,	5'd10,	5'd2};
		rom[ 1987 ] = { 5'd1,	5'd21,	5'd10,	5'd2};
		rom[ 1988 ] = { 5'd6,	5'd20,	5'd18,	5'd1};
		rom[ 1989 ] = { 5'd8,	5'd19,	5'd4,	5'd5};
		rom[ 1990 ] = { 5'd0,	5'd2,	5'd24,	5'd2};
		rom[ 1991 ] = { 5'd0,	5'd4,	5'd6,	5'd3};
		rom[ 1992 ] = { 5'd14,	5'd9,	5'd10,	5'd3};
		rom[ 1993 ] = { 5'd1,	5'd19,	5'd19,	5'd4};
		rom[ 1994 ] = { 5'd14,	5'd2,	5'd10,	5'd2};
		rom[ 1995 ] = { 5'd8,	5'd10,	5'd7,	5'd14};
		rom[ 1996 ] = { 5'd10,	5'd10,	5'd4,	5'd8};
		rom[ 1997 ] = { 5'd11,	5'd8,	5'd5,	5'd4};
		rom[ 1998 ] = { 5'd10,	5'd5,	5'd2,	5'd9};
		rom[ 1999 ] = { 5'd9,	5'd5,	5'd2,	5'd10};
		rom[ 2000 ] = { 5'd14,	5'd4,	5'd2,	5'd13};
		rom[ 2001 ] = { 5'd8,	5'd4,	5'd2,	5'd13};
		rom[ 2002 ] = { 5'd11,	5'd7,	5'd3,	5'd6};
		rom[ 2003 ] = { 5'd3,	5'd6,	5'd8,	5'd3};
		rom[ 2004 ] = { 5'd13,	5'd4,	5'd8,	5'd7};
		rom[ 2005 ] = { 5'd0,	5'd0,	5'd12,	5'd2};
		rom[ 2006 ] = { 5'd12,	5'd1,	5'd3,	5'd6};
		rom[ 2007 ] = { 5'd11,	5'd1,	5'd7,	5'd4};
		rom[ 2008 ] = { 5'd10,	5'd17,	5'd7,	5'd3};
		rom[ 2009 ] = { 5'd8,	5'd3,	5'd4,	5'd5};
		rom[ 2010 ] = { 5'd11,	5'd3,	5'd4,	5'd5};
		rom[ 2011 ] = { 5'd10,	5'd2,	5'd2,	5'd13};
		rom[ 2012 ] = { 5'd12,	5'd2,	5'd1,	5'd19};
		rom[ 2013 ] = { 5'd10,	5'd7,	5'd3,	5'd6};
		rom[ 2014 ] = { 5'd4,	5'd22,	5'd10,	5'd2};
		rom[ 2015 ] = { 5'd0,	5'd16,	5'd12,	5'd2};
		rom[ 2016 ] = { 5'd11,	5'd3,	5'd4,	5'd5};
		rom[ 2017 ] = { 5'd1,	5'd10,	5'd4,	5'd7};
		rom[ 2018 ] = { 5'd11,	5'd19,	5'd6,	5'd3};
		rom[ 2019 ] = { 5'd6,	5'd0,	5'd5,	5'd12};
		rom[ 2020 ] = { 5'd14,	5'd5,	5'd7,	5'd7};
		rom[ 2021 ] = { 5'd7,	5'd8,	5'd5,	5'd4};
		rom[ 2022 ] = { 5'd12,	5'd1,	5'd3,	5'd6};
		rom[ 2023 ] = { 5'd12,	5'd6,	5'd12,	5'd3};
		rom[ 2024 ] = { 5'd11,	5'd3,	5'd4,	5'd5};
		rom[ 2025 ] = { 5'd1,	5'd13,	5'd11,	5'd2};
		rom[ 2026 ] = { 5'd9,	5'd14,	5'd12,	5'd2};
		rom[ 2027 ] = { 5'd0,	5'd7,	5'd9,	5'd2};
		rom[ 2028 ] = { 5'd1,	5'd7,	5'd23,	5'd2};
		rom[ 2029 ] = { 5'd1,	5'd10,	5'd19,	5'd4};
		rom[ 2030 ] = { 5'd9,	5'd8,	5'd6,	5'd7};
		rom[ 2031 ] = { 5'd9,	5'd19,	5'd6,	5'd3};
		rom[ 2032 ] = { 5'd11,	5'd14,	5'd2,	5'd9};
		rom[ 2033 ] = { 5'd11,	5'd6,	5'd2,	5'd12};
		rom[ 2034 ] = { 5'd18,	5'd0,	5'd2,	5'd9};
		rom[ 2035 ] = { 5'd4,	5'd0,	5'd2,	5'd9};
		rom[ 2036 ] = { 5'd15,	5'd1,	5'd2,	5'd11};
		rom[ 2037 ] = { 5'd1,	5'd14,	5'd8,	5'd6};
		rom[ 2038 ] = { 5'd14,	5'd10,	5'd7,	5'd3};
		rom[ 2039 ] = { 5'd3,	5'd12,	5'd9,	5'd2};
		rom[ 2040 ] = { 5'd15,	5'd1,	5'd2,	5'd11};
		rom[ 2041 ] = { 5'd7,	5'd1,	5'd2,	5'd11};
		rom[ 2042 ] = { 5'd14,	5'd7,	5'd10,	5'd2};
		rom[ 2043 ] = { 5'd12,	5'd10,	5'd3,	5'd7};
		rom[ 2044 ] = { 5'd7,	5'd7,	5'd5,	5'd4};
		rom[ 2045 ] = { 5'd0,	5'd8,	5'd4,	5'd5};
		rom[ 2046 ] = { 5'd19,	5'd0,	5'd4,	5'd6};
		rom[ 2047 ] = { 5'd1,	5'd0,	5'd4,	5'd6};
		rom[ 2048 ] = { 5'd16,	5'd5,	5'd2,	5'd16};
		rom[ 2049 ] = { 5'd6,	5'd5,	5'd2,	5'd16};
		rom[ 2050 ] = { 5'd17,	5'd0,	5'd2,	5'd16};
		rom[ 2051 ] = { 5'd5,	5'd0,	5'd2,	5'd16};
		rom[ 2052 ] = { 5'd0,	5'd3,	5'd24,	5'd1};
		rom[ 2053 ] = { 5'd7,	5'd3,	5'd10,	5'd2};
		rom[ 2054 ] = { 5'd1,	5'd4,	5'd23,	5'd4};
		rom[ 2055 ] = { 5'd1,	5'd18,	5'd19,	5'd1};
		rom[ 2056 ] = { 5'd6,	5'd19,	5'd18,	5'd1};
		rom[ 2057 ] = { 5'd1,	5'd19,	5'd9,	5'd2};
		rom[ 2058 ] = { 5'd15,	5'd18,	5'd6,	5'd3};
		rom[ 2059 ] = { 5'd3,	5'd18,	5'd6,	5'd3};
		rom[ 2060 ] = { 5'd4,	5'd17,	5'd20,	5'd3};
		rom[ 2061 ] = { 5'd0,	5'd10,	5'd3,	5'd7};
		rom[ 2062 ] = { 5'd6,	5'd19,	5'd18,	5'd1};
		rom[ 2063 ] = { 5'd7,	5'd12,	5'd3,	5'd7};
		rom[ 2064 ] = { 5'd12,	5'd10,	5'd6,	5'd5};
		rom[ 2065 ] = { 5'd6,	5'd10,	5'd6,	5'd5};
		rom[ 2066 ] = { 5'd9,	5'd2,	5'd6,	5'd9};
		rom[ 2067 ] = { 5'd4,	5'd6,	5'd5,	5'd5};
		rom[ 2068 ] = { 5'd20,	5'd14,	5'd2,	5'd9};
		rom[ 2069 ] = { 5'd2,	5'd14,	5'd2,	5'd9};
		rom[ 2070 ] = { 5'd13,	5'd1,	5'd2,	5'd10};
		rom[ 2071 ] = { 5'd12,	5'd21,	5'd6,	5'd3};
		rom[ 2072 ] = { 5'd13,	5'd1,	5'd2,	5'd10};
		rom[ 2073 ] = { 5'd1,	5'd16,	5'd5,	5'd4};
		rom[ 2074 ] = { 5'd13,	5'd1,	5'd2,	5'd10};
		rom[ 2075 ] = { 5'd2,	5'd0,	5'd1,	5'd19};
		rom[ 2076 ] = { 5'd13,	5'd1,	5'd2,	5'd10};
		rom[ 2077 ] = { 5'd2,	5'd1,	5'd2,	5'd9};
		rom[ 2078 ] = { 5'd3,	5'd9,	5'd19,	5'd2};
		rom[ 2079 ] = { 5'd7,	5'd16,	5'd9,	5'd2};
		rom[ 2080 ] = { 5'd17,	5'd4,	5'd7,	5'd3};
		rom[ 2081 ] = { 5'd5,	5'd4,	5'd14,	5'd4};
		rom[ 2082 ] = { 5'd16,	5'd4,	5'd8,	5'd3};
		rom[ 2083 ] = { 5'd0,	5'd4,	5'd8,	5'd3};
		rom[ 2084 ] = { 5'd15,	5'd0,	5'd9,	5'd2};
		rom[ 2085 ] = { 5'd0,	5'd16,	5'd9,	5'd2};
		rom[ 2086 ] = { 5'd9,	5'd7,	5'd6,	5'd8};
		rom[ 2087 ] = { 5'd4,	5'd11,	5'd2,	5'd9};
		rom[ 2088 ] = { 5'd12,	5'd5,	5'd2,	5'd9};
		rom[ 2089 ] = { 5'd10,	5'd6,	5'd2,	5'd9};
		rom[ 2090 ] = { 5'd13,	5'd1,	5'd2,	5'd10};
		rom[ 2091 ] = { 5'd9,	5'd1,	5'd2,	5'd10};
		rom[ 2092 ] = { 5'd14,	5'd9,	5'd9,	5'd3};
		rom[ 2093 ] = { 5'd8,	5'd4,	5'd2,	5'd9};
		rom[ 2094 ] = { 5'd10,	5'd16,	5'd4,	5'd6};
		rom[ 2095 ] = { 5'd0,	5'd0,	5'd9,	5'd4};
		rom[ 2096 ] = { 5'd13,	5'd5,	5'd7,	5'd6};
		rom[ 2097 ] = { 5'd9,	5'd3,	5'd5,	5'd7};
		rom[ 2098 ] = { 5'd14,	5'd14,	5'd10,	5'd2};
		rom[ 2099 ] = { 5'd0,	5'd16,	5'd4,	5'd5};
		rom[ 2100 ] = { 5'd1,	5'd11,	5'd22,	5'd1};
		rom[ 2101 ] = { 5'd10,	5'd9,	5'd2,	5'd10};
		rom[ 2102 ] = { 5'd16,	5'd2,	5'd3,	5'd6};
		rom[ 2103 ] = { 5'd10,	5'd6,	5'd2,	5'd9};
		rom[ 2104 ] = { 5'd12,	5'd8,	5'd5,	5'd8};
		rom[ 2105 ] = { 5'd8,	5'd1,	5'd4,	5'd6};
		rom[ 2106 ] = { 5'd13,	5'd1,	5'd6,	5'd7};
		rom[ 2107 ] = { 5'd2,	5'd16,	5'd12,	5'd2};
		rom[ 2108 ] = { 5'd11,	5'd19,	5'd6,	5'd3};
		rom[ 2109 ] = { 5'd7,	5'd19,	5'd6,	5'd3};
		rom[ 2110 ] = { 5'd13,	5'd4,	5'd2,	5'd10};
		rom[ 2111 ] = { 5'd0,	5'd20,	5'd19,	5'd1};
		rom[ 2112 ] = { 5'd12,	5'd12,	5'd6,	5'd4};
		rom[ 2113 ] = { 5'd8,	5'd12,	5'd8,	5'd11};
		rom[ 2114 ] = { 5'd12,	5'd12,	5'd6,	5'd4};
		rom[ 2115 ] = { 5'd6,	5'd12,	5'd6,	5'd4};
		rom[ 2116 ] = { 5'd14,	5'd8,	5'd6,	5'd3};
		rom[ 2117 ] = { 5'd0,	5'd8,	5'd24,	5'd2};
		rom[ 2118 ] = { 5'd14,	5'd14,	5'd10,	5'd2};
		rom[ 2119 ] = { 5'd0,	5'd14,	5'd10,	5'd2};
		rom[ 2120 ] = { 5'd4,	5'd7,	5'd19,	5'd1};
		rom[ 2121 ] = { 5'd1,	5'd7,	5'd19,	5'd1};
		rom[ 2122 ] = { 5'd4,	5'd3,	5'd16,	5'd3};
		rom[ 2123 ] = { 5'd8,	5'd1,	5'd8,	5'd5};
		rom[ 2124 ] = { 5'd3,	5'd11,	5'd6,	5'd5};
		rom[ 2125 ] = { 5'd11,	5'd6,	5'd2,	5'd9};
		rom[ 2126 ] = { 5'd0,	5'd18,	5'd18,	5'd1};
		rom[ 2127 ] = { 5'd6,	5'd23,	5'd18,	5'd1};
		rom[ 2128 ] = { 5'd2,	5'd15,	5'd6,	5'd3};
		rom[ 2129 ] = { 5'd18,	5'd15,	5'd6,	5'd3};
		rom[ 2130 ] = { 5'd0,	5'd15,	5'd6,	5'd3};
		rom[ 2131 ] = { 5'd11,	5'd19,	5'd4,	5'd5};
		rom[ 2132 ] = { 5'd9,	5'd14,	5'd6,	5'd8};
		rom[ 2133 ] = { 5'd7,	5'd12,	5'd10,	5'd5};
		rom[ 2134 ] = { 5'd3,	5'd3,	5'd2,	5'd13};
		rom[ 2135 ] = { 5'd18,	5'd1,	5'd3,	5'd13};
		rom[ 2136 ] = { 5'd7,	5'd1,	5'd2,	5'd9};
		rom[ 2137 ] = { 5'd18,	5'd2,	5'd3,	5'd11};
		rom[ 2138 ] = { 5'd3,	5'd2,	5'd3,	5'd11};
		rom[ 2139 ] = { 5'd9,	5'd14,	5'd15,	5'd2};
		rom[ 2140 ] = { 5'd2,	5'd3,	5'd20,	5'd1};
		rom[ 2141 ] = { 5'd10,	5'd6,	5'd2,	5'd9};
		rom[ 2142 ] = { 5'd5,	5'd6,	5'd6,	5'd7};
		rom[ 2143 ] = { 5'd11,	5'd0,	5'd2,	5'd9};
		rom[ 2144 ] = { 5'd10,	5'd0,	5'd3,	5'd6};
		rom[ 2145 ] = { 5'd12,	5'd6,	5'd2,	5'd9};
		rom[ 2146 ] = { 5'd4,	5'd1,	5'd6,	5'd10};
		rom[ 2147 ] = { 5'd6,	5'd7,	5'd9,	5'd3};
		rom[ 2148 ] = { 5'd9,	5'd7,	5'd9,	5'd3};
		rom[ 2149 ] = { 5'd9,	5'd20,	5'd6,	5'd3};
		rom[ 2150 ] = { 5'd11,	5'd6,	5'd2,	5'd9};
		rom[ 2151 ] = { 5'd10,	5'd2,	5'd4,	5'd15};
		rom[ 2152 ] = { 5'd2,	5'd4,	5'd18,	5'd1};
		rom[ 2153 ] = { 5'd21,	5'd4,	5'd2,	5'd9};
		rom[ 2154 ] = { 5'd0,	5'd2,	5'd19,	5'd1};
		rom[ 2155 ] = { 5'd5,	5'd2,	5'd15,	5'd2};
		rom[ 2156 ] = { 5'd12,	5'd2,	5'd7,	5'd5};
		rom[ 2157 ] = { 5'd1,	5'd2,	5'd11,	5'd14};
		rom[ 2158 ] = { 5'd10,	5'd15,	5'd2,	5'd9};
		rom[ 2159 ] = { 5'd6,	5'd18,	5'd18,	5'd1};
		rom[ 2160 ] = { 5'd9,	5'd12,	5'd3,	5'd6};
		rom[ 2161 ] = { 5'd2,	5'd1,	5'd20,	5'd1};
		rom[ 2162 ] = { 5'd5,	5'd8,	5'd5,	5'd4};
		rom[ 2163 ] = { 5'd12,	5'd6,	5'd4,	5'd5};
		rom[ 2164 ] = { 5'd9,	5'd12,	5'd3,	5'd6};
		rom[ 2165 ] = { 5'd18,	5'd14,	5'd4,	5'd5};
		rom[ 2166 ] = { 5'd2,	5'd14,	5'd4,	5'd5};
		rom[ 2167 ] = { 5'd16,	5'd18,	5'd6,	5'd3};
		rom[ 2168 ] = { 5'd1,	5'd6,	5'd6,	5'd3};
		rom[ 2169 ] = { 5'd12,	5'd3,	5'd1,	5'd20};
		rom[ 2170 ] = { 5'd4,	5'd6,	5'd7,	5'd3};
		rom[ 2171 ] = { 5'd10,	5'd5,	5'd4,	5'd13};
		rom[ 2172 ] = { 5'd5,	5'd9,	5'd4,	5'd5};
		rom[ 2173 ] = { 5'd14,	5'd16,	5'd5,	5'd4};
		rom[ 2174 ] = { 5'd7,	5'd8,	5'd3,	5'd7};
		rom[ 2175 ] = { 5'd7,	5'd8,	5'd10,	5'd2};
		rom[ 2176 ] = { 5'd2,	5'd6,	5'd18,	5'd1};
		rom[ 2177 ] = { 5'd5,	5'd5,	5'd15,	5'd4};
		rom[ 2178 ] = { 5'd7,	5'd10,	5'd8,	5'd9};
		rom[ 2179 ] = { 5'd0,	5'd11,	5'd24,	5'd1};
		rom[ 2180 ] = { 5'd2,	5'd2,	5'd2,	5'd13};
		rom[ 2181 ] = { 5'd20,	5'd0,	5'd4,	5'd5};
		rom[ 2182 ] = { 5'd5,	5'd4,	5'd10,	5'd3};
		rom[ 2183 ] = { 5'd5,	5'd7,	5'd18,	5'd1};
		rom[ 2184 ] = { 5'd0,	5'd2,	5'd24,	5'd1};
		rom[ 2185 ] = { 5'd13,	5'd4,	5'd2,	5'd11};
		rom[ 2186 ] = { 5'd0,	5'd0,	5'd4,	5'd5};
		rom[ 2187 ] = { 5'd4,	5'd17,	5'd18,	5'd1};
		rom[ 2188 ] = { 5'd2,	5'd17,	5'd18,	5'd1};
		rom[ 2189 ] = { 5'd12,	5'd0,	5'd9,	5'd5};
		rom[ 2190 ] = { 5'd12,	5'd3,	5'd10,	5'd21};
		rom[ 2191 ] = { 5'd6,	5'd7,	5'd7,	5'd3};
		rom[ 2192 ] = { 5'd0,	5'd9,	5'd6,	5'd3};
		rom[ 2193 ] = { 5'd10,	5'd14,	5'd7,	5'd4};
		rom[ 2194 ] = { 5'd7,	5'd14,	5'd7,	5'd4};
		rom[ 2195 ] = { 5'd11,	5'd21,	5'd6,	5'd3};
		rom[ 2196 ] = { 5'd7,	5'd21,	5'd6,	5'd3};
		rom[ 2197 ] = { 5'd21,	5'd4,	5'd2,	5'd9};
		rom[ 2198 ] = { 5'd3,	5'd8,	5'd18,	5'd1};
		rom[ 2199 ] = { 5'd21,	5'd4,	5'd2,	5'd9};
		rom[ 2200 ] = { 5'd7,	5'd17,	5'd10,	5'd2};
		rom[ 2201 ] = { 5'd9,	5'd16,	5'd11,	5'd3};
		rom[ 2202 ] = { 5'd0,	5'd11,	5'd4,	5'd5};
		rom[ 2203 ] = { 5'd15,	5'd18,	5'd9,	5'd2};
		rom[ 2204 ] = { 5'd1,	5'd5,	5'd2,	5'd9};
		rom[ 2205 ] = { 5'd13,	5'd8,	5'd4,	5'd5};
		rom[ 2206 ] = { 5'd7,	5'd8,	5'd4,	5'd5};
		rom[ 2207 ] = { 5'd13,	5'd8,	5'd4,	5'd5};
		rom[ 2208 ] = { 5'd10,	5'd8,	5'd3,	5'd7};
		rom[ 2209 ] = { 5'd13,	5'd8,	5'd4,	5'd5};
		rom[ 2210 ] = { 5'd10,	5'd6,	5'd3,	5'd7};
		rom[ 2211 ] = { 5'd13,	5'd8,	5'd4,	5'd5};
		rom[ 2212 ] = { 5'd10,	5'd11,	5'd4,	5'd6};
		rom[ 2213 ] = { 5'd5,	5'd11,	5'd14,	5'd6};
		rom[ 2214 ] = { 5'd0,	5'd3,	5'd11,	5'd2};
		rom[ 2215 ] = { 5'd11,	5'd10,	5'd2,	5'd10};
		rom[ 2216 ] = { 5'd2,	5'd19,	5'd11,	5'd2};
		rom[ 2217 ] = { 5'd15,	5'd18,	5'd9,	5'd2};
		rom[ 2218 ] = { 5'd1,	5'd11,	5'd18,	5'd1};
		rom[ 2219 ] = { 5'd10,	5'd4,	5'd4,	5'd13};
		rom[ 2220 ] = { 5'd0,	5'd19,	5'd18,	5'd1};
		rom[ 2221 ] = { 5'd6,	5'd19,	5'd18,	5'd1};
		rom[ 2222 ] = { 5'd0,	5'd18,	5'd9,	5'd2};
		rom[ 2223 ] = { 5'd13,	5'd17,	5'd9,	5'd2};
		rom[ 2224 ] = { 5'd2,	5'd17,	5'd9,	5'd2};
		rom[ 2225 ] = { 5'd13,	5'd1,	5'd3,	5'd16};
		rom[ 2226 ] = { 5'd8,	5'd1,	5'd3,	5'd16};
		rom[ 2227 ] = { 5'd13,	5'd5,	5'd2,	5'd10};
		rom[ 2228 ] = { 5'd9,	5'd5,	5'd2,	5'd10};
		rom[ 2229 ] = { 5'd12,	5'd0,	5'd2,	5'd24};
		rom[ 2230 ] = { 5'd3,	5'd4,	5'd2,	5'd10};
		rom[ 2231 ] = { 5'd16,	5'd0,	5'd2,	5'd9};
		rom[ 2232 ] = { 5'd6,	5'd0,	5'd2,	5'd9};
		rom[ 2233 ] = { 5'd10,	5'd5,	5'd6,	5'd5};
		rom[ 2234 ] = { 5'd7,	5'd6,	5'd2,	5'd9};
		rom[ 2235 ] = { 5'd12,	5'd2,	5'd5,	5'd8};
		rom[ 2236 ] = { 5'd7,	5'd2,	5'd5,	5'd8};
		rom[ 2237 ] = { 5'd10,	5'd0,	5'd2,	5'd9};
		rom[ 2238 ] = { 5'd3,	5'd4,	5'd3,	5'd6};
		rom[ 2239 ] = { 5'd16,	5'd0,	5'd4,	5'd18};
		rom[ 2240 ] = { 5'd4,	5'd0,	5'd4,	5'd18};
		rom[ 2241 ] = { 5'd0,	5'd9,	5'd24,	5'd2};
		rom[ 2242 ] = { 5'd11,	5'd7,	5'd7,	5'd3};
		rom[ 2243 ] = { 5'd10,	5'd8,	5'd4,	5'd15};
		rom[ 2244 ] = { 5'd12,	5'd0,	5'd5,	5'd14};
		rom[ 2245 ] = { 5'd17,	5'd10,	5'd4,	5'd5};
		rom[ 2246 ] = { 5'd5,	5'd0,	5'd2,	5'd9};
		rom[ 2247 ] = { 5'd16,	5'd1,	5'd3,	5'd8};
		rom[ 2248 ] = { 5'd5,	5'd1,	5'd3,	5'd8};
		rom[ 2249 ] = { 5'd3,	5'd10,	5'd18,	5'd4};
		rom[ 2250 ] = { 5'd4,	5'd14,	5'd16,	5'd2};
		rom[ 2251 ] = { 5'd4,	5'd14,	5'd16,	5'd5};
		rom[ 2252 ] = { 5'd3,	5'd10,	5'd4,	5'd5};
		rom[ 2253 ] = { 5'd16,	5'd18,	5'd8,	5'd3};
		rom[ 2254 ] = { 5'd6,	5'd16,	5'd4,	5'd5};
		rom[ 2255 ] = { 5'd14,	5'd16,	5'd9,	5'd2};
		rom[ 2256 ] = { 5'd7,	5'd16,	5'd9,	5'd2};
		rom[ 2257 ] = { 5'd4,	5'd14,	5'd16,	5'd4};
		rom[ 2258 ] = { 5'd0,	5'd15,	5'd19,	5'd2};
		rom[ 2259 ] = { 5'd10,	5'd15,	5'd9,	5'd2};
		rom[ 2260 ] = { 5'd6,	5'd0,	5'd1,	5'd23};
		rom[ 2261 ] = { 5'd0,	5'd10,	5'd24,	5'd2};
		rom[ 2262 ] = { 5'd0,	5'd9,	5'd5,	5'd4};
		rom[ 2263 ] = { 5'd3,	5'd9,	5'd19,	5'd9};
		rom[ 2264 ] = { 5'd9,	5'd11,	5'd3,	5'd6};
		rom[ 2265 ] = { 5'd12,	5'd5,	5'd12,	5'd4};
		rom[ 2266 ] = { 5'd6,	5'd20,	5'd9,	5'd2};
		rom[ 2267 ] = { 5'd8,	5'd10,	5'd10,	5'd2};
		rom[ 2268 ] = { 5'd2,	5'd8,	5'd20,	5'd1};
		rom[ 2269 ] = { 5'd12,	5'd10,	5'd7,	5'd10};
		rom[ 2270 ] = { 5'd5,	5'd10,	5'd7,	5'd10};
		rom[ 2271 ] = { 5'd14,	5'd11,	5'd2,	5'd9};
		rom[ 2272 ] = { 5'd10,	5'd8,	5'd5,	5'd12};
		rom[ 2273 ] = { 5'd12,	5'd9,	5'd6,	5'd4};
		rom[ 2274 ] = { 5'd7,	5'd14,	5'd3,	5'd7};
		rom[ 2275 ] = { 5'd17,	5'd2,	5'd6,	5'd8};
		rom[ 2276 ] = { 5'd9,	5'd0,	5'd2,	5'd9};
		rom[ 2277 ] = { 5'd13,	5'd16,	5'd9,	5'd2};
		rom[ 2278 ] = { 5'd0,	5'd12,	5'd11,	5'd2};
		rom[ 2279 ] = { 5'd12,	5'd12,	5'd11,	5'd3};
		rom[ 2280 ] = { 5'd9,	5'd6,	5'd3,	5'd6};
		rom[ 2281 ] = { 5'd10,	5'd0,	5'd2,	5'd9};
		rom[ 2282 ] = { 5'd9,	5'd8,	5'd6,	5'd7};
		rom[ 2283 ] = { 5'd0,	5'd8,	5'd24,	5'd2};
		rom[ 2284 ] = { 5'd8,	5'd11,	5'd8,	5'd10};
		rom[ 2285 ] = { 5'd9,	5'd3,	5'd6,	5'd21};
		rom[ 2286 ] = { 5'd9,	5'd12,	5'd2,	5'd10};
		rom[ 2287 ] = { 5'd15,	5'd16,	5'd5,	5'd4};
		rom[ 2288 ] = { 5'd10,	5'd6,	5'd2,	5'd9};
		rom[ 2289 ] = { 5'd15,	5'd10,	5'd3,	5'd6};
		rom[ 2290 ] = { 5'd6,	5'd10,	5'd3,	5'd6};
		rom[ 2291 ] = { 5'd19,	5'd12,	5'd3,	5'd6};
		rom[ 2292 ] = { 5'd2,	5'd12,	5'd3,	5'd6};
		rom[ 2293 ] = { 5'd12,	5'd15,	5'd2,	5'd9};
		rom[ 2294 ] = { 5'd10,	5'd15,	5'd2,	5'd9};
		rom[ 2295 ] = { 5'd14,	5'd20,	5'd5,	5'd4};
		rom[ 2296 ] = { 5'd5,	5'd20,	5'd5,	5'd4};
		rom[ 2297 ] = { 5'd11,	5'd19,	5'd9,	5'd2};
		rom[ 2298 ] = { 5'd3,	5'd4,	5'd14,	5'd2};
		rom[ 2299 ] = { 5'd10,	5'd3,	5'd10,	5'd2};
		rom[ 2300 ] = { 5'd5,	5'd15,	5'd5,	5'd4};
		rom[ 2301 ] = { 5'd20,	5'd2,	5'd1,	5'd19};
		rom[ 2302 ] = { 5'd7,	5'd12,	5'd3,	5'd8};
		rom[ 2303 ] = { 5'd4,	5'd11,	5'd5,	5'd4};
		rom[ 2304 ] = { 5'd8,	5'd1,	5'd8,	5'd3};
		rom[ 2305 ] = { 5'd6,	5'd10,	5'd12,	5'd2};
		rom[ 2306 ] = { 5'd19,	5'd3,	5'd2,	5'd10};
		rom[ 2307 ] = { 5'd3,	5'd6,	5'd3,	5'd6};
		rom[ 2308 ] = { 5'd20,	5'd0,	5'd2,	5'd22};
		rom[ 2309 ] = { 5'd2,	5'd0,	5'd2,	5'd22};
		rom[ 2310 ] = { 5'd5,	5'd16,	5'd19,	5'd1};
		rom[ 2311 ] = { 5'd10,	5'd12,	5'd4,	5'd5};
		rom[ 2312 ] = { 5'd11,	5'd6,	5'd2,	5'd9};
		rom[ 2313 ] = { 5'd0,	5'd22,	5'd18,	5'd1};
		rom[ 2314 ] = { 5'd7,	5'd8,	5'd10,	5'd5};
		rom[ 2315 ] = { 5'd1,	5'd8,	5'd18,	5'd1};
		rom[ 2316 ] = { 5'd11,	5'd2,	5'd3,	5'd6};
		rom[ 2317 ] = { 5'd0,	5'd17,	5'd24,	5'd7};
		rom[ 2318 ] = { 5'd17,	5'd9,	5'd4,	5'd5};
		rom[ 2319 ] = { 5'd12,	5'd5,	5'd2,	5'd9};
		rom[ 2320 ] = { 5'd17,	5'd9,	5'd4,	5'd5};
		rom[ 2321 ] = { 5'd7,	5'd11,	5'd5,	5'd5};
		rom[ 2322 ] = { 5'd13,	5'd13,	5'd9,	5'd2};
		rom[ 2323 ] = { 5'd0,	5'd1,	5'd19,	5'd1};
		rom[ 2324 ] = { 5'd8,	5'd18,	5'd8,	5'd6};
		rom[ 2325 ] = { 5'd6,	5'd12,	5'd8,	5'd8};
		rom[ 2326 ] = { 5'd7,	5'd10,	5'd10,	5'd2};
		rom[ 2327 ] = { 5'd0,	5'd6,	5'd6,	5'd3};
		rom[ 2328 ] = { 5'd13,	5'd18,	5'd7,	5'd3};
		rom[ 2329 ] = { 5'd3,	5'd18,	5'd6,	5'd3};
		rom[ 2330 ] = { 5'd12,	5'd17,	5'd6,	5'd3};
		rom[ 2331 ] = { 5'd2,	5'd19,	5'd15,	5'd4};
		rom[ 2332 ] = { 5'd9,	5'd14,	5'd6,	5'd8};
		rom[ 2333 ] = { 5'd6,	5'd10,	5'd7,	5'd4};
		rom[ 2334 ] = { 5'd14,	5'd9,	5'd6,	5'd3};
		rom[ 2335 ] = { 5'd5,	5'd17,	5'd6,	5'd3};
		rom[ 2336 ] = { 5'd12,	5'd8,	5'd2,	5'd9};
		rom[ 2337 ] = { 5'd6,	5'd6,	5'd2,	5'd9};
		rom[ 2338 ] = { 5'd17,	5'd9,	5'd3,	5'd6};
		rom[ 2339 ] = { 5'd4,	5'd9,	5'd3,	5'd6};
		rom[ 2340 ] = { 5'd14,	5'd17,	5'd9,	5'd2};
		rom[ 2341 ] = { 5'd0,	5'd20,	5'd9,	5'd2};
		rom[ 2342 ] = { 5'd13,	5'd20,	5'd9,	5'd2};
		rom[ 2343 ] = { 5'd2,	5'd20,	5'd9,	5'd2};
		rom[ 2344 ] = { 5'd6,	5'd17,	5'd18,	5'd1};
		rom[ 2345 ] = { 5'd0,	5'd17,	5'd18,	5'd1};
		rom[ 2346 ] = { 5'd21,	5'd2,	5'd2,	5'd11};
		rom[ 2347 ] = { 5'd1,	5'd2,	5'd2,	5'd11};
		rom[ 2348 ] = { 5'd15,	5'd0,	5'd1,	5'd24};
		rom[ 2349 ] = { 5'd11,	5'd20,	5'd8,	5'd4};
		rom[ 2350 ] = { 5'd13,	5'd6,	5'd2,	5'd9};
		rom[ 2351 ] = { 5'd7,	5'd9,	5'd5,	5'd7};
		rom[ 2352 ] = { 5'd14,	5'd9,	5'd6,	5'd3};
		rom[ 2353 ] = { 5'd3,	5'd9,	5'd7,	5'd3};
		rom[ 2354 ] = { 5'd22,	5'd4,	5'd2,	5'd10};
		rom[ 2355 ] = { 5'd7,	5'd9,	5'd6,	5'd3};
		rom[ 2356 ] = { 5'd12,	5'd0,	5'd5,	5'd7};
		rom[ 2357 ] = { 5'd11,	5'd1,	5'd9,	5'd6};
		rom[ 2358 ] = { 5'd15,	5'd0,	5'd1,	5'd24};
		rom[ 2359 ] = { 5'd8,	5'd0,	5'd1,	5'd24};
		rom[ 2360 ] = { 5'd13,	5'd12,	5'd3,	5'd7};
		rom[ 2361 ] = { 5'd8,	5'd12,	5'd3,	5'd7};
		rom[ 2362 ] = { 5'd9,	5'd5,	5'd6,	5'd19};
		rom[ 2363 ] = { 5'd8,	5'd6,	5'd3,	5'd6};
		rom[ 2364 ] = { 5'd12,	5'd5,	5'd3,	5'd6};
		rom[ 2365 ] = { 5'd3,	5'd16,	5'd5,	5'd4};
		rom[ 2366 ] = { 5'd19,	5'd13,	5'd5,	5'd5};
		rom[ 2367 ] = { 5'd0,	5'd13,	5'd5,	5'd5};
		rom[ 2368 ] = { 5'd22,	5'd4,	5'd2,	5'd10};
		rom[ 2369 ] = { 5'd0,	5'd4,	5'd2,	5'd10};
		rom[ 2370 ] = { 5'd7,	5'd7,	5'd5,	5'd4};
		rom[ 2371 ] = { 5'd11,	5'd19,	5'd7,	5'd4};
		rom[ 2372 ] = { 5'd10,	5'd11,	5'd6,	5'd3};
		rom[ 2373 ] = { 5'd0,	5'd2,	5'd24,	5'd1};
		rom[ 2374 ] = { 5'd14,	5'd2,	5'd7,	5'd10};
		rom[ 2375 ] = { 5'd2,	5'd13,	5'd2,	5'd9};
		rom[ 2376 ] = { 5'd13,	5'd0,	5'd2,	5'd19};
		rom[ 2377 ] = { 5'd8,	5'd11,	5'd7,	5'd3};
		rom[ 2378 ] = { 5'd15,	5'd1,	5'd8,	5'd10};
		rom[ 2379 ] = { 5'd7,	5'd10,	5'd7,	5'd9};
		rom[ 2380 ] = { 5'd11,	5'd19,	5'd5,	5'd5};
		rom[ 2381 ] = { 5'd11,	5'd10,	5'd3,	5'd6};
		rom[ 2382 ] = { 5'd15,	5'd1,	5'd8,	5'd10};
		rom[ 2383 ] = { 5'd1,	5'd1,	5'd8,	5'd10};
		rom[ 2384 ] = { 5'd16,	5'd10,	5'd3,	5'd6};
		rom[ 2385 ] = { 5'd5,	5'd10,	5'd3,	5'd6};
		rom[ 2386 ] = { 5'd12,	5'd6,	5'd5,	5'd4};
		rom[ 2387 ] = { 5'd4,	5'd12,	5'd6,	5'd3};
		rom[ 2388 ] = { 5'd6,	5'd7,	5'd12,	5'd2};
		rom[ 2389 ] = { 5'd9,	5'd7,	5'd5,	5'd5};
		rom[ 2390 ] = { 5'd15,	5'd2,	5'd9,	5'd2};
		rom[ 2391 ] = { 5'd6,	5'd5,	5'd11,	5'd5};
		rom[ 2392 ] = { 5'd12,	5'd13,	5'd4,	5'd6};
		rom[ 2393 ] = { 5'd7,	5'd4,	5'd9,	5'd2};
		rom[ 2394 ] = { 5'd6,	5'd2,	5'd13,	5'd2};
		rom[ 2395 ] = { 5'd10,	5'd6,	5'd2,	5'd9};
		rom[ 2396 ] = { 5'd12,	5'd8,	5'd2,	5'd9};
		rom[ 2397 ] = { 5'd3,	5'd20,	5'd10,	5'd2};
		rom[ 2398 ] = { 5'd4,	5'd15,	5'd20,	5'd1};
		rom[ 2399 ] = { 5'd2,	5'd17,	5'd9,	5'd2};
		rom[ 2400 ] = { 5'd13,	5'd0,	5'd2,	5'd19};
		rom[ 2401 ] = { 5'd9,	5'd0,	5'd2,	5'd19};
		rom[ 2402 ] = { 5'd1,	5'd5,	5'd22,	5'd1};
		rom[ 2403 ] = { 5'd0,	5'd2,	5'd9,	5'd2};
		rom[ 2404 ] = { 5'd0,	5'd9,	5'd24,	5'd9};
		rom[ 2405 ] = { 5'd3,	5'd6,	5'd16,	5'd4};
		rom[ 2406 ] = { 5'd3,	5'd8,	5'd18,	5'd2};
		rom[ 2407 ] = { 5'd5,	5'd1,	5'd2,	5'd10};
		rom[ 2408 ] = { 5'd16,	5'd0,	5'd3,	5'd6};
		rom[ 2409 ] = { 5'd5,	5'd0,	5'd3,	5'd6};
		rom[ 2410 ] = { 5'd10,	5'd7,	5'd4,	5'd5};
		rom[ 2411 ] = { 5'd6,	5'd5,	5'd7,	5'd5};
		rom[ 2412 ] = { 5'd12,	5'd2,	5'd10,	5'd2};
		rom[ 2413 ] = { 5'd2,	5'd12,	5'd19,	5'd1};
		rom[ 2414 ] = { 5'd12,	5'd8,	5'd2,	5'd9};
		rom[ 2415 ] = { 5'd10,	5'd8,	5'd2,	5'd9};
		rom[ 2416 ] = { 5'd13,	5'd8,	5'd2,	5'd9};
		rom[ 2417 ] = { 5'd6,	5'd11,	5'd3,	5'd9};
		rom[ 2418 ] = { 5'd9,	5'd9,	5'd6,	5'd5};
		rom[ 2419 ] = { 5'd2,	5'd14,	5'd2,	5'd10};
		rom[ 2420 ] = { 5'd14,	5'd20,	5'd8,	5'd3};
		rom[ 2421 ] = { 5'd3,	5'd22,	5'd18,	5'd1};
		rom[ 2422 ] = { 5'd10,	5'd4,	5'd5,	5'd6};
		rom[ 2423 ] = { 5'd2,	5'd17,	5'd12,	5'd2};
		rom[ 2424 ] = { 5'd17,	5'd11,	5'd6,	5'd3};
		rom[ 2425 ] = { 5'd2,	5'd12,	5'd10,	5'd2};
		rom[ 2426 ] = { 5'd0,	5'd19,	5'd24,	5'd2};
		rom[ 2427 ] = { 5'd7,	5'd18,	5'd9,	5'd2};
		rom[ 2428 ] = { 5'd17,	5'd1,	5'd2,	5'd11};
		rom[ 2429 ] = { 5'd5,	5'd1,	5'd2,	5'd11};
		rom[ 2430 ] = { 5'd11,	5'd16,	5'd8,	5'd3};
		rom[ 2431 ] = { 5'd8,	5'd1,	5'd2,	5'd9};
		rom[ 2432 ] = { 5'd11,	5'd10,	5'd3,	5'd6};
		rom[ 2433 ] = { 5'd5,	5'd8,	5'd6,	5'd3};
		rom[ 2434 ] = { 5'd15,	5'd11,	5'd5,	5'd4};
		rom[ 2435 ] = { 5'd4,	5'd11,	5'd5,	5'd4};
		rom[ 2436 ] = { 5'd15,	5'd6,	5'd3,	5'd6};
		rom[ 2437 ] = { 5'd6,	5'd6,	5'd3,	5'd6};
		rom[ 2438 ] = { 5'd12,	5'd9,	5'd7,	5'd4};
		rom[ 2439 ] = { 5'd9,	5'd8,	5'd3,	5'd7};
		rom[ 2440 ] = { 5'd12,	5'd10,	5'd6,	5'd4};
		rom[ 2441 ] = { 5'd4,	5'd5,	5'd2,	5'd9};
		rom[ 2442 ] = { 5'd4,	5'd12,	5'd16,	5'd6};
		rom[ 2443 ] = { 5'd5,	5'd14,	5'd7,	5'd10};
		rom[ 2444 ] = { 5'd14,	5'd14,	5'd8,	5'd6};
		rom[ 2445 ] = { 5'd9,	5'd10,	5'd3,	5'd7};
		rom[ 2446 ] = { 5'd12,	5'd5,	5'd3,	5'd6};
		rom[ 2447 ] = { 5'd10,	5'd4,	5'd1,	5'd18};
		rom[ 2448 ] = { 5'd12,	5'd4,	5'd11,	5'd7};
		rom[ 2449 ] = { 5'd2,	5'd8,	5'd18,	5'd1};
		rom[ 2450 ] = { 5'd12,	5'd10,	5'd6,	5'd4};
		rom[ 2451 ] = { 5'd9,	5'd5,	5'd3,	5'd7};
		rom[ 2452 ] = { 5'd12,	5'd13,	5'd4,	5'd6};
		rom[ 2453 ] = { 5'd8,	5'd13,	5'd4,	5'd6};
		rom[ 2454 ] = { 5'd7,	5'd13,	5'd10,	5'd11};
		rom[ 2455 ] = { 5'd1,	5'd1,	5'd1,	5'd20};
		rom[ 2456 ] = { 5'd13,	5'd13,	5'd9,	5'd2};
		rom[ 2457 ] = { 5'd2,	5'd13,	5'd9,	5'd2};
		rom[ 2458 ] = { 5'd15,	5'd17,	5'd9,	5'd2};
		rom[ 2459 ] = { 5'd0,	5'd17,	5'd9,	5'd2};
		rom[ 2460 ] = { 5'd15,	5'd0,	5'd9,	5'd12};
		rom[ 2461 ] = { 5'd6,	5'd10,	5'd6,	5'd4};
		rom[ 2462 ] = { 5'd8,	5'd9,	5'd10,	5'd2};
		rom[ 2463 ] = { 5'd1,	5'd9,	5'd9,	5'd3};
		rom[ 2464 ] = { 5'd6,	5'd7,	5'd18,	5'd1};
		rom[ 2465 ] = { 5'd10,	5'd7,	5'd3,	5'd8};
		rom[ 2466 ] = { 5'd12,	5'd12,	5'd2,	5'd12};
		rom[ 2467 ] = { 5'd3,	5'd15,	5'd18,	5'd1};
		rom[ 2468 ] = { 5'd18,	5'd17,	5'd3,	5'd7};
		rom[ 2469 ] = { 5'd1,	5'd14,	5'd10,	5'd2};
		rom[ 2470 ] = { 5'd18,	5'd17,	5'd3,	5'd7};
		rom[ 2471 ] = { 5'd11,	5'd3,	5'd1,	5'd19};
		rom[ 2472 ] = { 5'd18,	5'd17,	5'd3,	5'd7};
		rom[ 2473 ] = { 5'd6,	5'd4,	5'd11,	5'd3};
		rom[ 2474 ] = { 5'd18,	5'd17,	5'd3,	5'd7};
		rom[ 2475 ] = { 5'd6,	5'd8,	5'd11,	5'd3};
		rom[ 2476 ] = { 5'd16,	5'd7,	5'd4,	5'd5};
		rom[ 2477 ] = { 5'd12,	5'd4,	5'd10,	5'd19};
		rom[ 2478 ] = { 5'd9,	5'd1,	5'd7,	5'd6};
		rom[ 2479 ] = { 5'd6,	5'd5,	5'd6,	5'd7};
		rom[ 2480 ] = { 5'd11,	5'd0,	5'd2,	5'd9};
		rom[ 2481 ] = { 5'd6,	5'd11,	5'd4,	5'd5};
		rom[ 2482 ] = { 5'd16,	5'd7,	5'd4,	5'd5};
		rom[ 2483 ] = { 5'd4,	5'd7,	5'd4,	5'd5};
		rom[ 2484 ] = { 5'd18,	5'd17,	5'd3,	5'd7};
		rom[ 2485 ] = { 5'd8,	5'd6,	5'd4,	5'd5};
		rom[ 2486 ] = { 5'd18,	5'd15,	5'd3,	5'd9};
		rom[ 2487 ] = { 5'd3,	5'd15,	5'd3,	5'd9};
		rom[ 2488 ] = { 5'd15,	5'd10,	5'd3,	5'd7};
		rom[ 2489 ] = { 5'd6,	5'd10,	5'd3,	5'd7};
		rom[ 2490 ] = { 5'd18,	5'd15,	5'd5,	5'd4};
		rom[ 2491 ] = { 5'd0,	5'd1,	5'd3,	5'd6};
		rom[ 2492 ] = { 5'd13,	5'd0,	5'd3,	5'd6};
		rom[ 2493 ] = { 5'd7,	5'd0,	5'd5,	5'd6};
		rom[ 2494 ] = { 5'd4,	5'd1,	5'd8,	5'd8};
		rom[ 2495 ] = { 5'd0,	5'd22,	5'd19,	5'd1};
		rom[ 2496 ] = { 5'd15,	5'd9,	5'd9,	5'd2};
		rom[ 2497 ] = { 5'd3,	5'd6,	5'd9,	5'd2};
		rom[ 2498 ] = { 5'd9,	5'd6,	5'd6,	5'd5};
		rom[ 2499 ] = { 5'd8,	5'd9,	5'd3,	5'd6};
		rom[ 2500 ] = { 5'd5,	5'd4,	5'd14,	5'd3};
		rom[ 2501 ] = { 5'd3,	5'd0,	5'd4,	5'd10};
		rom[ 2502 ] = { 5'd5,	5'd3,	5'd7,	5'd3};
		rom[ 2503 ] = { 5'd10,	5'd6,	5'd4,	5'd5};
		rom[ 2504 ] = { 5'd4,	5'd1,	5'd4,	5'd14};
		rom[ 2505 ] = { 5'd2,	5'd14,	5'd22,	5'd2};
		rom[ 2506 ] = { 5'd8,	5'd20,	5'd6,	5'd3};
		rom[ 2507 ] = { 5'd18,	5'd1,	5'd3,	5'd7};
		rom[ 2508 ] = { 5'd3,	5'd0,	5'd3,	5'd6};
		rom[ 2509 ] = { 5'd4,	5'd12,	5'd17,	5'd6};
		rom[ 2510 ] = { 5'd6,	5'd0,	5'd6,	5'd3};
		rom[ 2511 ] = { 5'd13,	5'd7,	5'd9,	5'd2};
		rom[ 2512 ] = { 5'd4,	5'd14,	5'd10,	5'd2};
		rom[ 2513 ] = { 5'd12,	5'd9,	5'd5,	5'd6};
		rom[ 2514 ] = { 5'd8,	5'd1,	5'd8,	5'd3};
		rom[ 2515 ] = { 5'd13,	5'd11,	5'd3,	5'd6};
		rom[ 2516 ] = { 5'd8,	5'd11,	5'd3,	5'd6};
		rom[ 2517 ] = { 5'd3,	5'd11,	5'd19,	5'd1};
		rom[ 2518 ] = { 5'd0,	5'd5,	5'd6,	5'd3};
		rom[ 2519 ] = { 5'd14,	5'd18,	5'd10,	5'd2};
		rom[ 2520 ] = { 5'd0,	5'd18,	5'd10,	5'd2};
		rom[ 2521 ] = { 5'd14,	5'd15,	5'd9,	5'd2};
		rom[ 2522 ] = { 5'd0,	5'd17,	5'd18,	5'd1};
		rom[ 2523 ] = { 5'd6,	5'd17,	5'd18,	5'd1};
		rom[ 2524 ] = { 5'd0,	5'd20,	5'd9,	5'd2};
		rom[ 2525 ] = { 5'd14,	5'd15,	5'd9,	5'd2};
		rom[ 2526 ] = { 5'd8,	5'd2,	5'd2,	5'd9};
		rom[ 2527 ] = { 5'd15,	5'd8,	5'd2,	5'd12};
		rom[ 2528 ] = { 5'd8,	5'd17,	5'd8,	5'd4};
		rom[ 2529 ] = { 5'd10,	5'd20,	5'd6,	5'd3};
		rom[ 2530 ] = { 5'd7,	5'd8,	5'd2,	5'd12};
		rom[ 2531 ] = { 5'd7,	5'd7,	5'd6,	5'd3};
		rom[ 2532 ] = { 5'd12,	5'd6,	5'd2,	5'd9};
		rom[ 2533 ] = { 5'd11,	5'd20,	5'd6,	5'd3};
		rom[ 2534 ] = { 5'd7,	5'd20,	5'd6,	5'd3};
		rom[ 2535 ] = { 5'd21,	5'd1,	5'd3,	5'd10};
		rom[ 2536 ] = { 5'd0,	5'd1,	5'd3,	5'd10};
		rom[ 2537 ] = { 5'd15,	5'd3,	5'd2,	5'd9};
		rom[ 2538 ] = { 5'd0,	5'd6,	5'd6,	5'd4};
		rom[ 2539 ] = { 5'd18,	5'd9,	5'd6,	5'd3};
		rom[ 2540 ] = { 5'd7,	5'd3,	5'd2,	5'd9};
		rom[ 2541 ] = { 5'd16,	5'd0,	5'd2,	5'd9};
		rom[ 2542 ] = { 5'd0,	5'd9,	5'd6,	5'd3};
		rom[ 2543 ] = { 5'd18,	5'd4,	5'd4,	5'd10};
		rom[ 2544 ] = { 5'd2,	5'd4,	5'd4,	5'd10};
		rom[ 2545 ] = { 5'd14,	5'd15,	5'd9,	5'd2};
		rom[ 2546 ] = { 5'd1,	5'd15,	5'd9,	5'd2};
		rom[ 2547 ] = { 5'd9,	5'd15,	5'd6,	5'd3};
		rom[ 2548 ] = { 5'd5,	5'd15,	5'd9,	5'd2};
		rom[ 2549 ] = { 5'd5,	5'd1,	5'd18,	5'd1};
		rom[ 2550 ] = { 5'd11,	5'd2,	5'd3,	5'd7};
		rom[ 2551 ] = { 5'd12,	5'd1,	5'd3,	5'd6};
		rom[ 2552 ] = { 5'd9,	5'd1,	5'd3,	5'd6};
		rom[ 2553 ] = { 5'd12,	5'd6,	5'd7,	5'd3};
		rom[ 2554 ] = { 5'd10,	5'd2,	5'd2,	5'd13};
		rom[ 2555 ] = { 5'd12,	5'd11,	5'd6,	5'd3};
		rom[ 2556 ] = { 5'd9,	5'd1,	5'd6,	5'd15};
		rom[ 2557 ] = { 5'd13,	5'd0,	5'd3,	5'd7};
		rom[ 2558 ] = { 5'd3,	5'd6,	5'd16,	5'd3};
		rom[ 2559 ] = { 5'd12,	5'd7,	5'd3,	5'd6};
		rom[ 2560 ] = { 5'd9,	5'd7,	5'd2,	5'd9};
		rom[ 2561 ] = { 5'd13,	5'd0,	5'd2,	5'd24};
		rom[ 2562 ] = { 5'd9,	5'd0,	5'd2,	5'd24};
		rom[ 2563 ] = { 5'd11,	5'd13,	5'd5,	5'd4};
		rom[ 2564 ] = { 5'd7,	5'd17,	5'd9,	5'd2};
		rom[ 2565 ] = { 5'd5,	5'd9,	5'd18,	5'd2};
		rom[ 2566 ] = { 5'd8,	5'd13,	5'd5,	5'd4};
		rom[ 2567 ] = { 5'd4,	5'd19,	5'd17,	5'd2};
		rom[ 2568 ] = { 5'd0,	5'd3,	5'd9,	5'd7};
		rom[ 2569 ] = { 5'd0,	5'd2,	5'd24,	5'd1};
		rom[ 2570 ] = { 5'd0,	5'd16,	5'd18,	5'd1};
		rom[ 2571 ] = { 5'd11,	5'd0,	5'd2,	5'd9};
		rom[ 2572 ] = { 5'd3,	5'd9,	5'd14,	5'd6};
		rom[ 2573 ] = { 5'd12,	5'd7,	5'd3,	5'd6};
		rom[ 2574 ] = { 5'd10,	5'd0,	5'd2,	5'd9};
		rom[ 2575 ] = { 5'd12,	5'd6,	5'd2,	5'd10};
		rom[ 2576 ] = { 5'd7,	5'd0,	5'd2,	5'd9};
		rom[ 2577 ] = { 5'd9,	5'd0,	5'd7,	5'd7};
		rom[ 2578 ] = { 5'd10,	5'd11,	5'd4,	5'd5};
		rom[ 2579 ] = { 5'd11,	5'd7,	5'd3,	5'd8};
		rom[ 2580 ] = { 5'd9,	5'd6,	5'd3,	5'd9};
		rom[ 2581 ] = { 5'd19,	5'd14,	5'd4,	5'd5};
		rom[ 2582 ] = { 5'd1,	5'd14,	5'd4,	5'd5};
		rom[ 2583 ] = { 5'd15,	5'd0,	5'd4,	5'd5};
		rom[ 2584 ] = { 5'd5,	5'd0,	5'd4,	5'd5};
		rom[ 2585 ] = { 5'd6,	5'd1,	5'd6,	5'd5};
		rom[ 2586 ] = { 5'd10,	5'd12,	5'd9,	5'd2};
		rom[ 2587 ] = { 5'd12,	5'd8,	5'd10,	5'd3};
		rom[ 2588 ] = { 5'd10,	5'd6,	5'd3,	5'd7};
		rom[ 2589 ] = { 5'd14,	5'd5,	5'd4,	5'd8};
		rom[ 2590 ] = { 5'd3,	5'd9,	5'd8,	5'd4};
		rom[ 2591 ] = { 5'd7,	5'd8,	5'd5,	5'd4};
		rom[ 2592 ] = { 5'd7,	5'd12,	5'd5,	5'd4};
		rom[ 2593 ] = { 5'd14,	5'd19,	5'd5,	5'd4};
		rom[ 2594 ] = { 5'd7,	5'd0,	5'd6,	5'd9};
		rom[ 2595 ] = { 5'd18,	5'd4,	5'd5,	5'd4};
		rom[ 2596 ] = { 5'd9,	5'd16,	5'd6,	5'd4};
		rom[ 2597 ] = { 5'd13,	5'd7,	5'd5,	5'd6};
		rom[ 2598 ] = { 5'd6,	5'd7,	5'd5,	5'd6};
		rom[ 2599 ] = { 5'd10,	5'd6,	5'd6,	5'd7};
		rom[ 2600 ] = { 5'd0,	5'd18,	5'd18,	5'd1};
		rom[ 2601 ] = { 5'd3,	5'd18,	5'd18,	5'd1};
		rom[ 2602 ] = { 5'd4,	5'd4,	5'd2,	5'd10};
		rom[ 2603 ] = { 5'd16,	5'd0,	5'd4,	5'd24};
		rom[ 2604 ] = { 5'd8,	5'd0,	5'd4,	5'd15};
		rom[ 2605 ] = { 5'd16,	5'd0,	5'd4,	5'd24};
		rom[ 2606 ] = { 5'd7,	5'd4,	5'd6,	5'd9};
		rom[ 2607 ] = { 5'd15,	5'd14,	5'd9,	5'd2};
		rom[ 2608 ] = { 5'd3,	5'd9,	5'd9,	5'd3};
		rom[ 2609 ] = { 5'd18,	5'd8,	5'd6,	5'd3};
		rom[ 2610 ] = { 5'd0,	5'd8,	5'd6,	5'd3};
		rom[ 2611 ] = { 5'd13,	5'd7,	5'd9,	5'd2};
		rom[ 2612 ] = { 5'd2,	5'd1,	5'd6,	5'd10};
		rom[ 2613 ] = { 5'd17,	5'd0,	5'd3,	5'd23};
		rom[ 2614 ] = { 5'd1,	5'd15,	5'd2,	5'd9};
		rom[ 2615 ] = { 5'd8,	5'd10,	5'd10,	5'd2};
		rom[ 2616 ] = { 5'd0,	5'd6,	5'd10,	5'd3};
		rom[ 2617 ] = { 5'd15,	5'd12,	5'd4,	5'd5};
		rom[ 2618 ] = { 5'd1,	5'd4,	5'd1,	5'd19};
		rom[ 2619 ] = { 5'd20,	5'd1,	5'd1,	5'd18};
		rom[ 2620 ] = { 5'd3,	5'd1,	5'd1,	5'd18};
		rom[ 2621 ] = { 5'd9,	5'd10,	5'd6,	5'd3};
		rom[ 2622 ] = { 5'd9,	5'd4,	5'd5,	5'd9};
		rom[ 2623 ] = { 5'd7,	5'd13,	5'd7,	5'd7};
		rom[ 2624 ] = { 5'd10,	5'd13,	5'd7,	5'd7};
		rom[ 2625 ] = { 5'd11,	5'd15,	5'd3,	5'd6};
		rom[ 2626 ] = { 5'd4,	5'd14,	5'd4,	5'd5};
		rom[ 2627 ] = { 5'd10,	5'd19,	5'd4,	5'd5};
		rom[ 2628 ] = { 5'd3,	5'd16,	5'd5,	5'd8};
		rom[ 2629 ] = { 5'd15,	5'd12,	5'd9,	5'd2};
		rom[ 2630 ] = { 5'd0,	5'd12,	5'd9,	5'd2};
		rom[ 2631 ] = { 5'd6,	5'd10,	5'd12,	5'd3};
		rom[ 2632 ] = { 5'd9,	5'd14,	5'd5,	5'd4};
		rom[ 2633 ] = { 5'd12,	5'd7,	5'd3,	5'd6};
		rom[ 2634 ] = { 5'd10,	5'd15,	5'd2,	5'd9};
		rom[ 2635 ] = { 5'd16,	5'd9,	5'd7,	5'd3};
		rom[ 2636 ] = { 5'd10,	5'd1,	5'd2,	5'd22};
		rom[ 2637 ] = { 5'd6,	5'd6,	5'd7,	5'd3};
		rom[ 2638 ] = { 5'd0,	5'd19,	5'd19,	5'd1};
		rom[ 2639 ] = { 5'd17,	5'd0,	5'd3,	5'd24};
		rom[ 2640 ] = { 5'd5,	5'd13,	5'd5,	5'd6};
		rom[ 2641 ] = { 5'd14,	5'd6,	5'd5,	5'd7};
		rom[ 2642 ] = { 5'd1,	5'd6,	5'd4,	5'd5};
		rom[ 2643 ] = { 5'd7,	5'd6,	5'd6,	5'd5};
		rom[ 2644 ] = { 5'd10,	5'd7,	5'd3,	5'd6};
		rom[ 2645 ] = { 5'd14,	5'd8,	5'd7,	5'd7};
		rom[ 2646 ] = { 5'd3,	5'd8,	5'd7,	5'd7};
		rom[ 2647 ] = { 5'd9,	5'd10,	5'd13,	5'd2};
		rom[ 2648 ] = { 5'd3,	5'd2,	5'd3,	5'd6};
		rom[ 2649 ] = { 5'd6,	5'd13,	5'd17,	5'd3};
		rom[ 2650 ] = { 5'd1,	5'd13,	5'd17,	5'd3};
		rom[ 2651 ] = { 5'd16,	5'd10,	5'd8,	5'd3};
		rom[ 2652 ] = { 5'd0,	5'd10,	5'd8,	5'd3};
		rom[ 2653 ] = { 5'd12,	5'd9,	5'd12,	5'd5};
		rom[ 2654 ] = { 5'd8,	5'd2,	5'd5,	5'd8};
		rom[ 2655 ] = { 5'd10,	5'd2,	5'd6,	5'd8};
		rom[ 2656 ] = { 5'd0,	5'd1,	5'd9,	5'd2};
		rom[ 2657 ] = { 5'd21,	5'd2,	5'd1,	5'd18};
		rom[ 2658 ] = { 5'd2,	5'd3,	5'd1,	5'd19};
		rom[ 2659 ] = { 5'd20,	5'd8,	5'd2,	5'd16};
		rom[ 2660 ] = { 5'd2,	5'd8,	5'd2,	5'd16};
		rom[ 2661 ] = { 5'd8,	5'd20,	5'd11,	5'd2};
		rom[ 2662 ] = { 5'd8,	5'd6,	5'd4,	5'd5};
		rom[ 2663 ] = { 5'd11,	5'd6,	5'd4,	5'd5};
		rom[ 2664 ] = { 5'd9,	5'd3,	5'd3,	5'd6};
		rom[ 2665 ] = { 5'd7,	5'd6,	5'd6,	5'd5};
		rom[ 2666 ] = { 5'd12,	5'd8,	5'd3,	5'd7};
		rom[ 2667 ] = { 5'd11,	5'd2,	5'd3,	5'd6};
		rom[ 2668 ] = { 5'd8,	5'd17,	5'd6,	5'd3};
		rom[ 2669 ] = { 5'd11,	5'd2,	5'd3,	5'd6};
		rom[ 2670 ] = { 5'd4,	5'd3,	5'd8,	5'd10};
		rom[ 2671 ] = { 5'd12,	5'd6,	5'd5,	5'd6};
		rom[ 2672 ] = { 5'd0,	5'd6,	5'd7,	5'd4};
		rom[ 2673 ] = { 5'd12,	5'd19,	5'd11,	5'd2};
		rom[ 2674 ] = { 5'd4,	5'd7,	5'd6,	5'd4};
		rom[ 2675 ] = { 5'd12,	5'd11,	5'd4,	5'd5};
		rom[ 2676 ] = { 5'd11,	5'd1,	5'd2,	5'd9};
		rom[ 2677 ] = { 5'd15,	5'd0,	5'd1,	5'd22};
		rom[ 2678 ] = { 5'd8,	5'd0,	5'd1,	5'd22};
		rom[ 2679 ] = { 5'd13,	5'd7,	5'd9,	5'd2};
		rom[ 2680 ] = { 5'd10,	5'd7,	5'd4,	5'd5};
		rom[ 2681 ] = { 5'd12,	5'd7,	5'd3,	5'd6};
		rom[ 2682 ] = { 5'd9,	5'd0,	5'd9,	5'd13};
		rom[ 2683 ] = { 5'd17,	5'd0,	5'd1,	5'd24};
		rom[ 2684 ] = { 5'd6,	5'd0,	5'd1,	5'd24};
		rom[ 2685 ] = { 5'd10,	5'd19,	5'd5,	5'd4};
		rom[ 2686 ] = { 5'd2,	5'd19,	5'd18,	5'd1};
		rom[ 2687 ] = { 5'd2,	5'd9,	5'd20,	5'd1};
		rom[ 2688 ] = { 5'd7,	5'd8,	5'd9,	5'd2};
		rom[ 2689 ] = { 5'd3,	5'd7,	5'd19,	5'd5};
		rom[ 2690 ] = { 5'd2,	5'd8,	5'd19,	5'd1};
		rom[ 2691 ] = { 5'd15,	5'd8,	5'd9,	5'd2};
		rom[ 2692 ] = { 5'd8,	5'd2,	5'd6,	5'd8};
		rom[ 2693 ] = { 5'd10,	5'd9,	5'd7,	5'd4};
		rom[ 2694 ] = { 5'd7,	5'd4,	5'd3,	5'd16};
		rom[ 2695 ] = { 5'd18,	5'd8,	5'd3,	5'd16};
		rom[ 2696 ] = { 5'd3,	5'd8,	5'd3,	5'd16};
		rom[ 2697 ] = { 5'd20,	5'd0,	5'd2,	5'd14};
		rom[ 2698 ] = { 5'd2,	5'd0,	5'd2,	5'd14};
		rom[ 2699 ] = { 5'd17,	5'd0,	5'd2,	5'd22};
		rom[ 2700 ] = { 5'd5,	5'd0,	5'd2,	5'd22};
		rom[ 2701 ] = { 5'd16,	5'd2,	5'd4,	5'd20};
		rom[ 2702 ] = { 5'd4,	5'd2,	5'd4,	5'd20};
		rom[ 2703 ] = { 5'd11,	5'd6,	5'd2,	5'd9};
		rom[ 2704 ] = { 5'd12,	5'd0,	5'd3,	5'd16};
		rom[ 2705 ] = { 5'd12,	5'd7,	5'd3,	5'd6};
		rom[ 2706 ] = { 5'd3,	5'd4,	5'd9,	5'd3};
		rom[ 2707 ] = { 5'd13,	5'd5,	5'd8,	5'd4};
		rom[ 2708 ] = { 5'd0,	5'd15,	5'd10,	5'd2};
		rom[ 2709 ] = { 5'd8,	5'd16,	5'd9,	5'd2};
		rom[ 2710 ] = { 5'd9,	5'd2,	5'd3,	5'd6};
		rom[ 2711 ] = { 5'd19,	5'd1,	5'd5,	5'd4};
		rom[ 2712 ] = { 5'd9,	5'd7,	5'd3,	5'd6};
		rom[ 2713 ] = { 5'd6,	5'd7,	5'd12,	5'd3};
		rom[ 2714 ] = { 5'd10,	5'd5,	5'd4,	5'd6};
		rom[ 2715 ] = { 5'd5,	5'd1,	5'd4,	5'd5};
		rom[ 2716 ] = { 5'd12,	5'd16,	5'd6,	5'd4};
		rom[ 2717 ] = { 5'd3,	5'd14,	5'd12,	5'd2};
		rom[ 2718 ] = { 5'd15,	5'd18,	5'd6,	5'd3};
		rom[ 2719 ] = { 5'd4,	5'd16,	5'd6,	5'd3};
		rom[ 2720 ] = { 5'd11,	5'd12,	5'd7,	5'd9};
		rom[ 2721 ] = { 5'd9,	5'd9,	5'd6,	5'd3};
		rom[ 2722 ] = { 5'd5,	5'd4,	5'd19,	5'd1};
		rom[ 2723 ] = { 5'd4,	5'd2,	5'd6,	5'd3};
		rom[ 2724 ] = { 5'd11,	5'd6,	5'd2,	5'd9};
		rom[ 2725 ] = { 5'd10,	5'd6,	5'd2,	5'd9};
		rom[ 2726 ] = { 5'd16,	5'd14,	5'd5,	5'd5};
		rom[ 2727 ] = { 5'd3,	5'd14,	5'd5,	5'd5};
		rom[ 2728 ] = { 5'd13,	5'd6,	5'd7,	5'd3};
		rom[ 2729 ] = { 5'd8,	5'd13,	5'd3,	5'd7};
		rom[ 2730 ] = { 5'd8,	5'd16,	5'd8,	5'd5};
		rom[ 2731 ] = { 5'd10,	5'd20,	5'd10,	5'd3};
		rom[ 2732 ] = { 5'd5,	5'd11,	5'd18,	5'd1};
		rom[ 2733 ] = { 5'd2,	5'd6,	5'd2,	5'd10};
		rom[ 2734 ] = { 5'd2,	5'd2,	5'd20,	5'd1};
		rom[ 2735 ] = { 5'd11,	5'd13,	5'd2,	5'd11};
		rom[ 2736 ] = { 5'd9,	5'd19,	5'd6,	5'd4};
		rom[ 2737 ] = { 5'd9,	5'd15,	5'd6,	5'd3};
		rom[ 2738 ] = { 5'd5,	5'd12,	5'd18,	5'd1};
		rom[ 2739 ] = { 5'd2,	5'd8,	5'd15,	5'd2};
		rom[ 2740 ] = { 5'd6,	5'd1,	5'd18,	5'd1};
		rom[ 2741 ] = { 5'd6,	5'd0,	5'd1,	5'd18};
		rom[ 2742 ] = { 5'd20,	5'd3,	5'd2,	5'd10};
		rom[ 2743 ] = { 5'd2,	5'd3,	5'd2,	5'd10};
		rom[ 2744 ] = { 5'd10,	5'd5,	5'd4,	5'd9};
		rom[ 2745 ] = { 5'd10,	5'd5,	5'd4,	5'd9};
		rom[ 2746 ] = { 5'd3,	5'd3,	5'd20,	5'd1};
		rom[ 2747 ] = { 5'd5,	5'd4,	5'd13,	5'd2};
		rom[ 2748 ] = { 5'd17,	5'd7,	5'd7,	5'd7};
		rom[ 2749 ] = { 5'd0,	5'd7,	5'd7,	5'd7};
		rom[ 2750 ] = { 5'd9,	5'd11,	5'd5,	5'd6};
		rom[ 2751 ] = { 5'd10,	5'd11,	5'd5,	5'd6};
		rom[ 2752 ] = { 5'd11,	5'd12,	5'd3,	5'd6};
		rom[ 2753 ] = { 5'd0,	5'd17,	5'd18,	5'd1};
		rom[ 2754 ] = { 5'd6,	5'd17,	5'd18,	5'd1};
		rom[ 2755 ] = { 5'd4,	5'd11,	5'd9,	5'd5};
		rom[ 2756 ] = { 5'd9,	5'd9,	5'd15,	5'd2};
		rom[ 2757 ] = { 5'd5,	5'd6,	5'd6,	5'd3};
		rom[ 2758 ] = { 5'd6,	5'd4,	5'd12,	5'd3};
		rom[ 2759 ] = { 5'd7,	5'd9,	5'd3,	5'd6};
		rom[ 2760 ] = { 5'd11,	5'd7,	5'd13,	5'd2};
		rom[ 2761 ] = { 5'd12,	5'd11,	5'd11,	5'd13};
		rom[ 2762 ] = { 5'd18,	5'd11,	5'd6,	5'd3};
		rom[ 2763 ] = { 5'd0,	5'd11,	5'd6,	5'd3};
		rom[ 2764 ] = { 5'd0,	5'd7,	5'd24,	5'd1};
		rom[ 2765 ] = { 5'd0,	5'd7,	5'd10,	5'd2};
		rom[ 2766 ] = { 5'd6,	5'd8,	5'd18,	5'd1};
		rom[ 2767 ] = { 5'd0,	5'd2,	5'd10,	5'd2};
		rom[ 2768 ] = { 5'd20,	5'd0,	5'd1,	5'd19};
		rom[ 2769 ] = { 5'd4,	5'd6,	5'd6,	5'd8};
		rom[ 2770 ] = { 5'd21,	5'd6,	5'd2,	5'd9};
		rom[ 2771 ] = { 5'd1,	5'd6,	5'd2,	5'd9};
		rom[ 2772 ] = { 5'd3,	5'd22,	5'd18,	5'd1};
		rom[ 2773 ] = { 5'd0,	5'd21,	5'd9,	5'd2};
		rom[ 2774 ] = { 5'd18,	5'd18,	5'd6,	5'd3};
		rom[ 2775 ] = { 5'd7,	5'd20,	5'd9,	5'd2};
		rom[ 2776 ] = { 5'd17,	5'd16,	5'd5,	5'd4};
		rom[ 2777 ] = { 5'd2,	5'd16,	5'd5,	5'd4};
		rom[ 2778 ] = { 5'd19,	5'd0,	5'd5,	5'd6};
		rom[ 2779 ] = { 5'd0,	5'd0,	5'd5,	5'd6};
		rom[ 2780 ] = { 5'd15,	5'd16,	5'd9,	5'd2};
		rom[ 2781 ] = { 5'd0,	5'd16,	5'd9,	5'd2};
		rom[ 2782 ] = { 5'd14,	5'd16,	5'd10,	5'd2};
		rom[ 2783 ] = { 5'd0,	5'd16,	5'd10,	5'd2};
		rom[ 2784 ] = { 5'd5,	5'd19,	5'd18,	5'd1};
		rom[ 2785 ] = { 5'd0,	5'd19,	5'd18,	5'd1};
		rom[ 2786 ] = { 5'd12,	5'd5,	5'd9,	5'd6};
		rom[ 2787 ] = { 5'd5,	5'd6,	5'd7,	5'd3};
		rom[ 2788 ] = { 5'd4,	5'd5,	5'd19,	5'd5};
		rom[ 2789 ] = { 5'd3,	5'd2,	5'd16,	5'd2};
		rom[ 2790 ] = { 5'd4,	5'd12,	5'd8,	5'd12};
		rom[ 2791 ] = { 5'd10,	5'd3,	5'd6,	5'd15};
		rom[ 2792 ] = { 5'd16,	5'd4,	5'd1,	5'd19};
		rom[ 2793 ] = { 5'd7,	5'd4,	5'd1,	5'd19};
		rom[ 2794 ] = { 5'd17,	5'd14,	5'd4,	5'd5};
		rom[ 2795 ] = { 5'd3,	5'd14,	5'd4,	5'd5};
		rom[ 2796 ] = { 5'd12,	5'd12,	5'd3,	5'd6};
		rom[ 2797 ] = { 5'd5,	5'd11,	5'd6,	5'd3};
		rom[ 2798 ] = { 5'd14,	5'd5,	5'd4,	5'd5};
		rom[ 2799 ] = { 5'd6,	5'd4,	5'd6,	5'd5};
		rom[ 2800 ] = { 5'd15,	5'd8,	5'd9,	5'd5};
		rom[ 2801 ] = { 5'd0,	5'd8,	5'd9,	5'd5};
		rom[ 2802 ] = { 5'd12,	5'd12,	5'd3,	5'd6};
		rom[ 2803 ] = { 5'd0,	5'd15,	5'd18,	5'd1};
		rom[ 2804 ] = { 5'd12,	5'd12,	5'd3,	5'd6};
		rom[ 2805 ] = { 5'd9,	5'd12,	5'd3,	5'd6};
		rom[ 2806 ] = { 5'd6,	5'd15,	5'd18,	5'd1};
		rom[ 2807 ] = { 5'd0,	5'd6,	5'd18,	5'd1};
		rom[ 2808 ] = { 5'd2,	5'd6,	5'd22,	5'd1};
		rom[ 2809 ] = { 5'd7,	5'd0,	5'd7,	5'd10};
		rom[ 2810 ] = { 5'd12,	5'd3,	5'd6,	5'd17};
		rom[ 2811 ] = { 5'd6,	5'd3,	5'd6,	5'd17};
		rom[ 2812 ] = { 5'd8,	5'd12,	5'd8,	5'd11};
		rom[ 2813 ] = { 5'd4,	5'd13,	5'd16,	5'd3};
		rom[ 2814 ] = { 5'd12,	5'd12,	5'd6,	5'd4};
		rom[ 2815 ] = { 5'd10,	5'd14,	5'd4,	5'd7};
		rom[ 2816 ] = { 5'd18,	5'd10,	5'd3,	5'd7};
		rom[ 2817 ] = { 5'd3,	5'd10,	5'd3,	5'd7};
		rom[ 2818 ] = { 5'd6,	5'd13,	5'd18,	5'd1};
		rom[ 2819 ] = { 5'd5,	5'd10,	5'd10,	5'd2};
		rom[ 2820 ] = { 5'd12,	5'd13,	5'd9,	5'd2};
		rom[ 2821 ] = { 5'd0,	5'd13,	5'd9,	5'd2};
		rom[ 2822 ] = { 5'd12,	5'd2,	5'd1,	5'd18};
		rom[ 2823 ] = { 5'd11,	5'd2,	5'd1,	5'd18};
		rom[ 2824 ] = { 5'd11,	5'd12,	5'd2,	5'd10};
		rom[ 2825 ] = { 5'd1,	5'd13,	5'd6,	5'd3};
		rom[ 2826 ] = { 5'd14,	5'd9,	5'd8,	5'd3};
		rom[ 2827 ] = { 5'd1,	5'd10,	5'd9,	5'd2};
		rom[ 2828 ] = { 5'd7,	5'd9,	5'd16,	5'd2};
		rom[ 2829 ] = { 5'd0,	5'd1,	5'd18,	5'd1};
		rom[ 2830 ] = { 5'd12,	5'd0,	5'd2,	5'd9};
		rom[ 2831 ] = { 5'd12,	5'd5,	5'd3,	5'd6};
		rom[ 2832 ] = { 5'd12,	5'd6,	5'd2,	5'd9};
		rom[ 2833 ] = { 5'd10,	5'd0,	5'd2,	5'd9};
		rom[ 2834 ] = { 5'd9,	5'd4,	5'd6,	5'd3};
		rom[ 2835 ] = { 5'd1,	5'd3,	5'd18,	5'd3};
		rom[ 2836 ] = { 5'd0,	5'd4,	5'd24,	5'd1};
		rom[ 2837 ] = { 5'd6,	5'd16,	5'd9,	5'd2};
		rom[ 2838 ] = { 5'd12,	5'd9,	5'd4,	5'd5};
		rom[ 2839 ] = { 5'd5,	5'd5,	5'd13,	5'd3};
		rom[ 2840 ] = { 5'd4,	5'd7,	5'd16,	5'd3};
		rom[ 2841 ] = { 5'd4,	5'd7,	5'd14,	5'd3};
		rom[ 2842 ] = { 5'd8,	5'd7,	5'd9,	5'd2};
		rom[ 2843 ] = { 5'd1,	5'd9,	5'd16,	5'd2};
		rom[ 2844 ] = { 5'd10,	5'd8,	5'd13,	5'd3};
		rom[ 2845 ] = { 5'd1,	5'd8,	5'd13,	5'd3};
		rom[ 2846 ] = { 5'd12,	5'd4,	5'd12,	5'd3};
		rom[ 2847 ] = { 5'd1,	5'd17,	5'd10,	5'd3};
		rom[ 2848 ] = { 5'd5,	5'd18,	5'd18,	5'd1};
		rom[ 2849 ] = { 5'd0,	5'd17,	5'd18,	5'd1};
		rom[ 2850 ] = { 5'd9,	5'd19,	5'd9,	5'd2};
		rom[ 2851 ] = { 5'd1,	5'd20,	5'd11,	5'd2};
		rom[ 2852 ] = { 5'd8,	5'd17,	5'd8,	5'd3};
		rom[ 2853 ] = { 5'd8,	5'd11,	5'd8,	5'd5};
		rom[ 2854 ] = { 5'd5,	5'd5,	5'd18,	5'd1};
		rom[ 2855 ] = { 5'd9,	5'd8,	5'd5,	5'd5};
		rom[ 2856 ] = { 5'd6,	5'd8,	5'd6,	5'd3};
		rom[ 2857 ] = { 5'd2,	5'd6,	5'd9,	5'd3};
		rom[ 2858 ] = { 5'd12,	5'd6,	5'd2,	5'd9};
		rom[ 2859 ] = { 5'd10,	5'd5,	5'd3,	5'd6};
		rom[ 2860 ] = { 5'd14,	5'd14,	5'd2,	5'd9};
		rom[ 2861 ] = { 5'd8,	5'd14,	5'd2,	5'd9};
		rom[ 2862 ] = { 5'd9,	5'd2,	5'd5,	5'd6};
		rom[ 2863 ] = { 5'd12,	5'd1,	5'd9,	5'd12};
		rom[ 2864 ] = { 5'd5,	5'd13,	5'd17,	5'd11};
		rom[ 2865 ] = { 5'd4,	5'd2,	5'd12,	5'd2};
		rom[ 2866 ] = { 5'd14,	5'd9,	5'd8,	5'd3};
		rom[ 2867 ] = { 5'd9,	5'd9,	5'd5,	5'd9};
		rom[ 2868 ] = { 5'd14,	5'd0,	5'd2,	5'd9};
		rom[ 2869 ] = { 5'd8,	5'd0,	5'd2,	5'd9};
		rom[ 2870 ] = { 5'd11,	5'd1,	5'd2,	5'd12};
		rom[ 2871 ] = { 5'd5,	5'd11,	5'd13,	5'd2};
		rom[ 2872 ] = { 5'd5,	5'd9,	5'd19,	5'd1};
		rom[ 2873 ] = { 5'd9,	5'd13,	5'd6,	5'd4};
		rom[ 2874 ] = { 5'd11,	5'd14,	5'd4,	5'd5};
		rom[ 2875 ] = { 5'd2,	5'd0,	5'd3,	5'd7};
		rom[ 2876 ] = { 5'd18,	5'd1,	5'd3,	5'd7};
		rom[ 2877 ] = { 5'd3,	5'd1,	5'd3,	5'd7};
		rom[ 2878 ] = { 5'd12,	5'd20,	5'd9,	5'd2};
		rom[ 2879 ] = { 5'd5,	5'd0,	5'd2,	5'd10};
		rom[ 2880 ] = { 5'd20,	5'd8,	5'd4,	5'd6};
		rom[ 2881 ] = { 5'd0,	5'd8,	5'd4,	5'd6};
		rom[ 2882 ] = { 5'd18,	5'd13,	5'd5,	5'd4};
		rom[ 2883 ] = { 5'd1,	5'd13,	5'd5,	5'd4};
		rom[ 2884 ] = { 5'd15,	5'd13,	5'd4,	5'd5};
		rom[ 2885 ] = { 5'd5,	5'd13,	5'd4,	5'd5};
		rom[ 2886 ] = { 5'd6,	5'd15,	5'd16,	5'd4};
		rom[ 2887 ] = { 5'd2,	5'd15,	5'd16,	5'd4};
		rom[ 2888 ] = { 5'd14,	5'd15,	5'd7,	5'd3};
		rom[ 2889 ] = { 5'd10,	5'd8,	5'd3,	5'd7};
		rom[ 2890 ] = { 5'd13,	5'd13,	5'd9,	5'd2};
		rom[ 2891 ] = { 5'd3,	5'd13,	5'd17,	5'd3};
		rom[ 2892 ] = { 5'd13,	5'd13,	5'd8,	5'd5};
		rom[ 2893 ] = { 5'd3,	5'd13,	5'd8,	5'd5};
		rom[ 2894 ] = { 5'd16,	5'd14,	5'd5,	5'd4};
		rom[ 2895 ] = { 5'd0,	5'd18,	5'd11,	5'd3};
		rom[ 2896 ] = { 5'd0,	5'd16,	5'd12,	5'd4};
		rom[ 2897 ] = { 5'd12,	5'd20,	5'd6,	5'd3};
		rom[ 2898 ] = { 5'd21,	5'd12,	5'd3,	5'd6};
		rom[ 2899 ] = { 5'd0,	5'd12,	5'd3,	5'd6};
		rom[ 2900 ] = { 5'd15,	5'd19,	5'd9,	5'd2};
		rom[ 2901 ] = { 5'd1,	5'd6,	5'd11,	5'd5};
		rom[ 2902 ] = { 5'd15,	5'd19,	5'd9,	5'd2};
		rom[ 2903 ] = { 5'd0,	5'd19,	5'd18,	5'd1};
		rom[ 2904 ] = { 5'd3,	5'd16,	5'd19,	5'd1};
		rom[ 2905 ] = { 5'd0,	5'd14,	5'd18,	5'd1};
		rom[ 2906 ] = { 5'd15,	5'd19,	5'd9,	5'd2};
		rom[ 2907 ] = { 5'd0,	5'd19,	5'd9,	5'd2};
		rom[ 2908 ] = { 5'd12,	5'd19,	5'd9,	5'd2};
		rom[ 2909 ] = { 5'd3,	5'd19,	5'd9,	5'd2};
		rom[ 2910 ] = { 5'd17,	5'd2,	5'd1,	5'd20};
		rom[ 2911 ] = { 5'd0,	5'd17,	5'd24,	5'd4};
		rom[ 2912 ] = { 5'd12,	5'd1,	5'd3,	5'd11};
	end
endmodule

module rect2_rom(
	input 				clk,
	input		[11:0]	addr,
	output reg	[19:0]	q    // x y w h 5bit*4
	);
	reg					[19:0]	rom [4095:0];
	always @(posedge clk) q <= rom[addr];
	initial begin
	rom[ 0    ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1    ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2    ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 3    ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 4    ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 5    ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 6    ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 7    ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 8    ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 9    ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 10   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 11   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 12   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 13   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 14   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 15   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 16   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 17   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 18   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 19   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 20   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 21   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 22   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 23   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 24   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 25   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 26   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 27   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 28   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 29   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 30   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 31   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 32   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 33   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 34   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 35   ] = { 5'd12,	5'd12,	5'd7,	5'd6};
	rom[ 36   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 37   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 38   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 39   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 40   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 41   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 42   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 43   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 44   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 45   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 46   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 47   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 48   ] = { 5'd5,	5'd12,	5'd7,	5'd7};
	rom[ 49   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 50   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 51   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 52   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 53   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 54   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 55   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 56   ] = { 5'd8,	5'd20,	5'd6,	5'd3};
	rom[ 57   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 58   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 59   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 60   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 61   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 62   ] = { 5'd11,	5'd15,	5'd8,	5'd3};
	rom[ 63   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 64   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 65   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 66   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 67   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 68   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 69   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 70   ] = { 5'd11,	5'd12,	5'd10,	5'd7};
	rom[ 71   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 72   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 73   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 74   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 75   ] = { 5'd11,	5'd11,	5'd4,	5'd5};
	rom[ 76   ] = { 5'd12,	5'd12,	5'd7,	5'd7};
	rom[ 77   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 78   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 79   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 80   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 81   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 82   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 83   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 84   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 85   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 86   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 87   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 88   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 89   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 90   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 91   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 92   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 93   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 94   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 95   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 96   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 97   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 98   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 99   ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 100  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 101  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 102  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 103  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 104  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 105  ] = { 5'd2,	5'd19,	5'd10,	5'd3};
	rom[ 106  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 107  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 108  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 109  ] = { 5'd11,	5'd11,	5'd6,	5'd3};
	rom[ 110  ] = { 5'd6,	5'd11,	5'd6,	5'd3};
	rom[ 111  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 112  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 113  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 114  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 115  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 116  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 117  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 118  ] = { 5'd11,	5'd15,	5'd9,	5'd6};
	rom[ 119  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 120  ] = { 5'd12,	5'd11,	5'd7,	5'd5};
	rom[ 121  ] = { 5'd9,	5'd11,	5'd5,	5'd6};
	rom[ 122  ] = { 5'd10,	5'd11,	5'd6,	5'd6};
	rom[ 123  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 124  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 125  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 126  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 127  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 128  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 129  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 130  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 131  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 132  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 133  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 134  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 135  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 136  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 137  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 138  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 139  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 140  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 141  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 142  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 143  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 144  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 145  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 146  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 147  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 148  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 149  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 150  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 151  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 152  ] = { 5'd9,	5'd11,	5'd4,	5'd5};
	rom[ 153  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 154  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 155  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 156  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 157  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 158  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 159  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 160  ] = { 5'd12,	5'd8,	5'd5,	5'd8};
	rom[ 161  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 162  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 163  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 164  ] = { 5'd11,	5'd3,	5'd10,	5'd2};
	rom[ 165  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 166  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 167  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 168  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 169  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 170  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 171  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 172  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 173  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 174  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 175  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 176  ] = { 5'd12,	5'd15,	5'd12,	5'd2};
	rom[ 177  ] = { 5'd2,	5'd10,	5'd11,	5'd6};
	rom[ 178  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 179  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 180  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 181  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 182  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 183  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 184  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 185  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 186  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 187  ] = { 5'd9,	5'd13,	5'd4,	5'd9};
	rom[ 188  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 189  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 190  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 191  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 192  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 193  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 194  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 195  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 196  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 197  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 198  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 199  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 200  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 201  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 202  ] = { 5'd6,	5'd11,	5'd7,	5'd6};
	rom[ 203  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 204  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 205  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 206  ] = { 5'd2,	5'd14,	5'd11,	5'd2};
	rom[ 207  ] = { 5'd11,	5'd14,	5'd11,	5'd2};
	rom[ 208  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 209  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 210  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 211  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 212  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 213  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 214  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 215  ] = { 5'd9,	5'd8,	5'd8,	5'd3};
	rom[ 216  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 217  ] = { 5'd12,	5'd11,	5'd12,	5'd7};
	rom[ 218  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 219  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 220  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 221  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 222  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 223  ] = { 5'd9,	5'd21,	5'd7,	5'd3};
	rom[ 224  ] = { 5'd3,	5'd20,	5'd9,	5'd2};
	rom[ 225  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 226  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 227  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 228  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 229  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 230  ] = { 5'd7,	5'd16,	5'd5,	5'd7};
	rom[ 231  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 232  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 233  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 234  ] = { 5'd3,	5'd18,	5'd9,	5'd2};
	rom[ 235  ] = { 5'd11,	5'd9,	5'd7,	5'd3};
	rom[ 236  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 237  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 238  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 239  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 240  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 241  ] = { 5'd12,	5'd5,	5'd12,	5'd3};
	rom[ 242  ] = { 5'd1,	5'd5,	5'd11,	5'd4};
	rom[ 243  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 244  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 245  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 246  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 247  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 248  ] = { 5'd17,	5'd16,	5'd3,	5'd8};
	rom[ 249  ] = { 5'd11,	5'd17,	5'd10,	5'd2};
	rom[ 250  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 251  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 252  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 253  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 254  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 255  ] = { 5'd9,	5'd19,	5'd6,	5'd5};
	rom[ 256  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 257  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 258  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 259  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 260  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 261  ] = { 5'd6,	5'd7,	5'd3,	5'd6};
	rom[ 262  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 263  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 264  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 265  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 266  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 267  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 268  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 269  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 270  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 271  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 272  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 273  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 274  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 275  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 276  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 277  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 278  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 279  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 280  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 281  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 282  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 283  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 284  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 285  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 286  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 287  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 288  ] = { 5'd7,	5'd15,	5'd5,	5'd6};
	rom[ 289  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 290  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 291  ] = { 5'd5,	5'd6,	5'd3,	5'd6};
	rom[ 292  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 293  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 294  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 295  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 296  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 297  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 298  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 299  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 300  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 301  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 302  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 303  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 304  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 305  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 306  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 307  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 308  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 309  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 310  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 311  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 312  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 313  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 314  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 315  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 316  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 317  ] = { 5'd11,	5'd11,	5'd10,	5'd8};
	rom[ 318  ] = { 5'd12,	5'd11,	5'd3,	5'd6};
	rom[ 319  ] = { 5'd12,	5'd10,	5'd11,	5'd8};
	rom[ 320  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 321  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 322  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 323  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 324  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 325  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 326  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 327  ] = { 5'd8,	5'd19,	5'd4,	5'd5};
	rom[ 328  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 329  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 330  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 331  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 332  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 333  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 334  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 335  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 336  ] = { 5'd18,	5'd15,	5'd3,	5'd9};
	rom[ 337  ] = { 5'd3,	5'd15,	5'd3,	5'd9};
	rom[ 338  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 339  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 340  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 341  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 342  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 343  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 344  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 345  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 346  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 347  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 348  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 349  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 350  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 351  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 352  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 353  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 354  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 355  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 356  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 357  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 358  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 359  ] = { 5'd12,	5'd15,	5'd11,	5'd2};
	rom[ 360  ] = { 5'd4,	5'd9,	5'd8,	5'd3};
	rom[ 361  ] = { 5'd10,	5'd11,	5'd9,	5'd11};
	rom[ 362  ] = { 5'd10,	5'd14,	5'd4,	5'd7};
	rom[ 363  ] = { 5'd3,	5'd14,	5'd3,	5'd10};
	rom[ 364  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 365  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 366  ] = { 5'd15,	5'd18,	5'd3,	5'd6};
	rom[ 367  ] = { 5'd6,	5'd18,	5'd3,	5'd6};
	rom[ 368  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 369  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 370  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 371  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 372  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 373  ] = { 5'd11,	5'd6,	5'd5,	5'd6};
	rom[ 374  ] = { 5'd17,	5'd7,	5'd3,	5'd6};
	rom[ 375  ] = { 5'd4,	5'd7,	5'd3,	5'd6};
	rom[ 376  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 377  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 378  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 379  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 380  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 381  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 382  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 383  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 384  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 385  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 386  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 387  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 388  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 389  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 390  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 391  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 392  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 393  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 394  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 395  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 396  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 397  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 398  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 399  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 400  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 401  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 402  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 403  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 404  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 405  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 406  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 407  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 408  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 409  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 410  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 411  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 412  ] = { 5'd9,	5'd21,	5'd6,	5'd3};
	rom[ 413  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 414  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 415  ] = { 5'd8,	5'd13,	5'd5,	5'd6};
	rom[ 416  ] = { 5'd11,	5'd13,	5'd5,	5'd6};
	rom[ 417  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 418  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 419  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 420  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 421  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 422  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 423  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 424  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 425  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 426  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 427  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 428  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 429  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 430  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 431  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 432  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 433  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 434  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 435  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 436  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 437  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 438  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 439  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 440  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 441  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 442  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 443  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 444  ] = { 5'd12,	5'd9,	5'd7,	5'd3};
	rom[ 445  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 446  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 447  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 448  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 449  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 450  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 451  ] = { 5'd1,	5'd5,	5'd11,	5'd3};
	rom[ 452  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 453  ] = { 5'd0,	5'd8,	5'd12,	5'd8};
	rom[ 454  ] = { 5'd12,	5'd15,	5'd9,	5'd2};
	rom[ 455  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 456  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 457  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 458  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 459  ] = { 5'd14,	5'd5,	5'd5,	5'd5};
	rom[ 460  ] = { 5'd5,	5'd5,	5'd5,	5'd5};
	rom[ 461  ] = { 5'd0,	5'd3,	5'd12,	5'd2};
	rom[ 462  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 463  ] = { 5'd5,	5'd18,	5'd8,	5'd3};
	rom[ 464  ] = { 5'd11,	5'd18,	5'd8,	5'd3};
	rom[ 465  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 466  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 467  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 468  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 469  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 470  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 471  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 472  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 473  ] = { 5'd16,	5'd14,	5'd3,	5'd7};
	rom[ 474  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 475  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 476  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 477  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 478  ] = { 5'd5,	5'd14,	5'd3,	5'd7};
	rom[ 479  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 480  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 481  ] = { 5'd12,	5'd9,	5'd5,	5'd7};
	rom[ 482  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 483  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 484  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 485  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 486  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 487  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 488  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 489  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 490  ] = { 5'd12,	5'd15,	5'd2,	5'd9};
	rom[ 491  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 492  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 493  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 494  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 495  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 496  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 497  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 498  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 499  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 500  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 501  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 502  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 503  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 504  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 505  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 506  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 507  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 508  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 509  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 510  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 511  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 512  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 513  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 514  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 515  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 516  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 517  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 518  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 519  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 520  ] = { 5'd4,	5'd5,	5'd8,	5'd5};
	rom[ 521  ] = { 5'd7,	5'd8,	5'd5,	5'd8};
	rom[ 522  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 523  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 524  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 525  ] = { 5'd11,	5'd14,	5'd6,	5'd3};
	rom[ 526  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 527  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 528  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 529  ] = { 5'd11,	5'd17,	5'd4,	5'd5};
	rom[ 530  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 531  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 532  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 533  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 534  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 535  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 536  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 537  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 538  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 539  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 540  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 541  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 542  ] = { 5'd0,	5'd15,	5'd12,	5'd2};
	rom[ 543  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 544  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 545  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 546  ] = { 5'd16,	5'd17,	5'd4,	5'd7};
	rom[ 547  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 548  ] = { 5'd16,	5'd17,	5'd4,	5'd7};
	rom[ 549  ] = { 5'd4,	5'd17,	5'd4,	5'd7};
	rom[ 550  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 551  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 552  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 553  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 554  ] = { 5'd5,	5'd9,	5'd8,	5'd4};
	rom[ 555  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 556  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 557  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 558  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 559  ] = { 5'd6,	5'd18,	5'd4,	5'd5};
	rom[ 560  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 561  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 562  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 563  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 564  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 565  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 566  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 567  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 568  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 569  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 570  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 571  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 572  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 573  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 574  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 575  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 576  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 577  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 578  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 579  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 580  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 581  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 582  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 583  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 584  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 585  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 586  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 587  ] = { 5'd11,	5'd13,	5'd5,	5'd6};
	rom[ 588  ] = { 5'd10,	5'd15,	5'd2,	5'd9};
	rom[ 589  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 590  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 591  ] = { 5'd7,	5'd19,	5'd4,	5'd5};
	rom[ 592  ] = { 5'd0,	5'd14,	5'd12,	5'd2};
	rom[ 593  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 594  ] = { 5'd12,	5'd20,	5'd5,	5'd4};
	rom[ 595  ] = { 5'd7,	5'd20,	5'd5,	5'd4};
	rom[ 596  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 597  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 598  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 599  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 600  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 601  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 602  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 603  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 604  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 605  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 606  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 607  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 608  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 609  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 610  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 611  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 612  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 613  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 614  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 615  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 616  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 617  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 618  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 619  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 620  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 621  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 622  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 623  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 624  ] = { 5'd12,	5'd9,	5'd6,	5'd3};
	rom[ 625  ] = { 5'd8,	5'd13,	5'd4,	5'd5};
	rom[ 626  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 627  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 628  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 629  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 630  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 631  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 632  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 633  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 634  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 635  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 636  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 637  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 638  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 639  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 640  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 641  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 642  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 643  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 644  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 645  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 646  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 647  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 648  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 649  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 650  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 651  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 652  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 653  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 654  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 655  ] = { 5'd13,	5'd9,	5'd4,	5'd5};
	rom[ 656  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 657  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 658  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 659  ] = { 5'd7,	5'd9,	5'd7,	5'd3};
	rom[ 660  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 661  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 662  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 663  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 664  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 665  ] = { 5'd14,	5'd9,	5'd3,	5'd7};
	rom[ 666  ] = { 5'd7,	5'd9,	5'd3,	5'd7};
	rom[ 667  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 668  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 669  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 670  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 671  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 672  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 673  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 674  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 675  ] = { 5'd12,	5'd8,	5'd6,	5'd3};
	rom[ 676  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 677  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 678  ] = { 5'd6,	5'd8,	5'd6,	5'd3};
	rom[ 679  ] = { 5'd14,	5'd19,	5'd4,	5'd5};
	rom[ 680  ] = { 5'd6,	5'd19,	5'd4,	5'd5};
	rom[ 681  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 682  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 683  ] = { 5'd5,	5'd9,	5'd8,	5'd3};
	rom[ 684  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 685  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 686  ] = { 5'd10,	5'd11,	5'd7,	5'd6};
	rom[ 687  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 688  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 689  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 690  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 691  ] = { 5'd20,	5'd11,	5'd2,	5'd9};
	rom[ 692  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 693  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 694  ] = { 5'd2,	5'd11,	5'd2,	5'd9};
	rom[ 695  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 696  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 697  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 698  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 699  ] = { 5'd7,	5'd6,	5'd6,	5'd6};
	rom[ 700  ] = { 5'd12,	5'd6,	5'd12,	5'd3};
	rom[ 701  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 702  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 703  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 704  ] = { 5'd11,	5'd9,	5'd9,	5'd4};
	rom[ 705  ] = { 5'd7,	5'd9,	5'd7,	5'd3};
	rom[ 706  ] = { 5'd10,	5'd9,	5'd7,	5'd3};
	rom[ 707  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 708  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 709  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 710  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 711  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 712  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 713  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 714  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 715  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 716  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 717  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 718  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 719  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 720  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 721  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 722  ] = { 5'd17,	5'd6,	5'd3,	5'd6};
	rom[ 723  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 724  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 725  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 726  ] = { 5'd10,	5'd13,	5'd6,	5'd3};
	rom[ 727  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 728  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 729  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 730  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 731  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 732  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 733  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 734  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 735  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 736  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 737  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 738  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 739  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 740  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 741  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 742  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 743  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 744  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 745  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 746  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 747  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 748  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 749  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 750  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 751  ] = { 5'd12,	5'd16,	5'd7,	5'd7};
	rom[ 752  ] = { 5'd0,	5'd5,	5'd12,	5'd5};
	rom[ 753  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 754  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 755  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 756  ] = { 5'd16,	5'd15,	5'd4,	5'd9};
	rom[ 757  ] = { 5'd4,	5'd15,	5'd4,	5'd9};
	rom[ 758  ] = { 5'd12,	5'd11,	5'd6,	5'd6};
	rom[ 759  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 760  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 761  ] = { 5'd6,	5'd11,	5'd6,	5'd6};
	rom[ 762  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 763  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 764  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 765  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 766  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 767  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 768  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 769  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 770  ] = { 5'd3,	5'd14,	5'd10,	5'd4};
	rom[ 771  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 772  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 773  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 774  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 775  ] = { 5'd12,	5'd7,	5'd5,	5'd7};
	rom[ 776  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 777  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 778  ] = { 5'd13,	5'd15,	5'd4,	5'd5};
	rom[ 779  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 780  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 781  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 782  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 783  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 784  ] = { 5'd0,	5'd6,	5'd12,	5'd3};
	rom[ 785  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 786  ] = { 5'd0,	5'd2,	5'd12,	5'd2};
	rom[ 787  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 788  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 789  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 790  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 791  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 792  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 793  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 794  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 795  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 796  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 797  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 798  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 799  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 800  ] = { 5'd13,	5'd12,	5'd5,	5'd4};
	rom[ 801  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 802  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 803  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 804  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 805  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 806  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 807  ] = { 5'd11,	5'd10,	5'd3,	5'd7};
	rom[ 808  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 809  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 810  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 811  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 812  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 813  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 814  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 815  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 816  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 817  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 818  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 819  ] = { 5'd7,	5'd15,	5'd4,	5'd5};
	rom[ 820  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 821  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 822  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 823  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 824  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 825  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 826  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 827  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 828  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 829  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 830  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 831  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 832  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 833  ] = { 5'd11,	5'd8,	5'd4,	5'd6};
	rom[ 834  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 835  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 836  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 837  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 838  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 839  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 840  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 841  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 842  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 843  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 844  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 845  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 846  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 847  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 848  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 849  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 850  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 851  ] = { 5'd0,	5'd3,	5'd12,	5'd2};
	rom[ 852  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 853  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 854  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 855  ] = { 5'd1,	5'd11,	5'd11,	5'd6};
	rom[ 856  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 857  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 858  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 859  ] = { 5'd6,	5'd15,	5'd8,	5'd3};
	rom[ 860  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 861  ] = { 5'd11,	5'd15,	5'd3,	5'd7};
	rom[ 862  ] = { 5'd10,	5'd15,	5'd8,	5'd3};
	rom[ 863  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 864  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 865  ] = { 5'd8,	5'd7,	5'd4,	5'd5};
	rom[ 866  ] = { 5'd12,	5'd9,	5'd6,	5'd3};
	rom[ 867  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 868  ] = { 5'd4,	5'd6,	5'd4,	5'd6};
	rom[ 869  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 870  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 871  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 872  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 873  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 874  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 875  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 876  ] = { 5'd10,	5'd15,	5'd3,	5'd7};
	rom[ 877  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 878  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 879  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 880  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 881  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 882  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 883  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 884  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 885  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 886  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 887  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 888  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 889  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 890  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 891  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 892  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 893  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 894  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 895  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 896  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 897  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 898  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 899  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 900  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 901  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 902  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 903  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 904  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 905  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 906  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 907  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 908  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 909  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 910  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 911  ] = { 5'd8,	5'd8,	5'd4,	5'd5};
	rom[ 912  ] = { 5'd11,	5'd9,	5'd8,	5'd3};
	rom[ 913  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 914  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 915  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 916  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 917  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 918  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 919  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 920  ] = { 5'd5,	5'd13,	5'd3,	5'd8};
	rom[ 921  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 922  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 923  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 924  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 925  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 926  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 927  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 928  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 929  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 930  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 931  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 932  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 933  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 934  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 935  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 936  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 937  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 938  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 939  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 940  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 941  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 942  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 943  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 944  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 945  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 946  ] = { 5'd12,	5'd15,	5'd7,	5'd7};
	rom[ 947  ] = { 5'd1,	5'd19,	5'd11,	5'd3};
	rom[ 948  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 949  ] = { 5'd9,	5'd10,	5'd5,	5'd5};
	rom[ 950  ] = { 5'd10,	5'd10,	5'd5,	5'd5};
	rom[ 951  ] = { 5'd4,	5'd9,	5'd8,	5'd3};
	rom[ 952  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 953  ] = { 5'd16,	5'd17,	5'd4,	5'd7};
	rom[ 954  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 955  ] = { 5'd8,	5'd16,	5'd4,	5'd6};
	rom[ 956  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 957  ] = { 5'd10,	5'd12,	5'd4,	5'd8};
	rom[ 958  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 959  ] = { 5'd5,	5'd13,	5'd7,	5'd7};
	rom[ 960  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 961  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 962  ] = { 5'd7,	5'd16,	5'd6,	5'd5};
	rom[ 963  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 964  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 965  ] = { 5'd10,	5'd12,	5'd4,	5'd8};
	rom[ 966  ] = { 5'd10,	5'd12,	5'd4,	5'd8};
	rom[ 967  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 968  ] = { 5'd9,	5'd11,	5'd8,	5'd6};
	rom[ 969  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 970  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 971  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 972  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 973  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 974  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 975  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 976  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 977  ] = { 5'd9,	5'd21,	5'd6,	5'd3};
	rom[ 978  ] = { 5'd16,	5'd16,	5'd4,	5'd8};
	rom[ 979  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 980  ] = { 5'd16,	5'd16,	5'd4,	5'd8};
	rom[ 981  ] = { 5'd4,	5'd16,	5'd4,	5'd8};
	rom[ 982  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 983  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 984  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 985  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 986  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 987  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 988  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 989  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 990  ] = { 5'd6,	5'd15,	5'd6,	5'd4};
	rom[ 991  ] = { 5'd6,	5'd11,	5'd6,	5'd3};
	rom[ 992  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 993  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 994  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 995  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 996  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 997  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 998  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 999  ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1000 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1001 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1002 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1003 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1004 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1005 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1006 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1007 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1008 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1009 ] = { 5'd11,	5'd9,	5'd6,	5'd4};
	rom[ 1010 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1011 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1012 ] = { 5'd8,	5'd7,	5'd4,	5'd6};
	rom[ 1013 ] = { 5'd4,	5'd6,	5'd3,	5'd6};
	rom[ 1014 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1015 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1016 ] = { 5'd17,	5'd17,	5'd3,	5'd7};
	rom[ 1017 ] = { 5'd4,	5'd17,	5'd3,	5'd7};
	rom[ 1018 ] = { 5'd7,	5'd13,	5'd7,	5'd7};
	rom[ 1019 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1020 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1021 ] = { 5'd12,	5'd3,	5'd11,	5'd2};
	rom[ 1022 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1023 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1024 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1025 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1026 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1027 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1028 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1029 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1030 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1031 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1032 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1033 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1034 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1035 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1036 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1037 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1038 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1039 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1040 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1041 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1042 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1043 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1044 ] = { 5'd3,	5'd15,	5'd9,	5'd2};
	rom[ 1045 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1046 ] = { 5'd4,	5'd3,	5'd10,	5'd2};
	rom[ 1047 ] = { 5'd10,	5'd3,	5'd10,	5'd2};
	rom[ 1048 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1049 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1050 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1051 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1052 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1053 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1054 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1055 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1056 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1057 ] = { 5'd11,	5'd16,	5'd4,	5'd7};
	rom[ 1058 ] = { 5'd1,	5'd8,	5'd11,	5'd3};
	rom[ 1059 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1060 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1061 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1062 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1063 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1064 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1065 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1066 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1067 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1068 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1069 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1070 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1071 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1072 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1073 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1074 ] = { 5'd12,	5'd14,	5'd5,	5'd4};
	rom[ 1075 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1076 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1077 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1078 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1079 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1080 ] = { 5'd9,	5'd14,	5'd7,	5'd5};
	rom[ 1081 ] = { 5'd8,	5'd14,	5'd7,	5'd5};
	rom[ 1082 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1083 ] = { 5'd6,	5'd14,	5'd3,	5'd10};
	rom[ 1084 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1085 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1086 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1087 ] = { 5'd6,	5'd16,	5'd3,	5'd8};
	rom[ 1088 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1089 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1090 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1091 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1092 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1093 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1094 ] = { 5'd12,	5'd20,	5'd5,	5'd4};
	rom[ 1095 ] = { 5'd7,	5'd20,	5'd5,	5'd4};
	rom[ 1096 ] = { 5'd0,	5'd2,	5'd12,	5'd2};
	rom[ 1097 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1098 ] = { 5'd0,	5'd7,	5'd12,	5'd3};
	rom[ 1099 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1100 ] = { 5'd1,	5'd3,	5'd11,	5'd2};
	rom[ 1101 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1102 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1103 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1104 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1105 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1106 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1107 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1108 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1109 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1110 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1111 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1112 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1113 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1114 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1115 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1116 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1117 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1118 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1119 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1120 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1121 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1122 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1123 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1124 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1125 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1126 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1127 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1128 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1129 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1130 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1131 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1132 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1133 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1134 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1135 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1136 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1137 ] = { 5'd12,	5'd12,	5'd7,	5'd7};
	rom[ 1138 ] = { 5'd12,	5'd11,	5'd6,	5'd3};
	rom[ 1139 ] = { 5'd12,	5'd12,	5'd6,	5'd6};
	rom[ 1140 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1141 ] = { 5'd11,	5'd14,	5'd10,	5'd4};
	rom[ 1142 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1143 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1144 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1145 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1146 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1147 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1148 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1149 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1150 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1151 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1152 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1153 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1154 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1155 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1156 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1157 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1158 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1159 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1160 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1161 ] = { 5'd12,	5'd4,	5'd11,	5'd2};
	rom[ 1162 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1163 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1164 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1165 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1166 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1167 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1168 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1169 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1170 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1171 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1172 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1173 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1174 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1175 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1176 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1177 ] = { 5'd12,	5'd11,	5'd12,	5'd8};
	rom[ 1178 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1179 ] = { 5'd11,	5'd9,	5'd6,	5'd4};
	rom[ 1180 ] = { 5'd5,	5'd9,	5'd7,	5'd3};
	rom[ 1181 ] = { 5'd12,	5'd19,	5'd7,	5'd3};
	rom[ 1182 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1183 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1184 ] = { 5'd3,	5'd9,	5'd10,	5'd5};
	rom[ 1185 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1186 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1187 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1188 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1189 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1190 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1191 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1192 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1193 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1194 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1195 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1196 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1197 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1198 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1199 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1200 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1201 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1202 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1203 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1204 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1205 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1206 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1207 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1208 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1209 ] = { 5'd8,	5'd21,	5'd8,	5'd3};
	rom[ 1210 ] = { 5'd9,	5'd21,	5'd7,	5'd3};
	rom[ 1211 ] = { 5'd11,	5'd22,	5'd10,	5'd2};
	rom[ 1212 ] = { 5'd2,	5'd11,	5'd10,	5'd3};
	rom[ 1213 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1214 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1215 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1216 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1217 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1218 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1219 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1220 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1221 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1222 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1223 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1224 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1225 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1226 ] = { 5'd10,	5'd5,	5'd4,	5'd5};
	rom[ 1227 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1228 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1229 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1230 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1231 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1232 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1233 ] = { 5'd6,	5'd5,	5'd6,	5'd5};
	rom[ 1234 ] = { 5'd10,	5'd4,	5'd6,	5'd3};
	rom[ 1235 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1236 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1237 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1238 ] = { 5'd6,	5'd5,	5'd6,	5'd3};
	rom[ 1239 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1240 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1241 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1242 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1243 ] = { 5'd4,	5'd18,	5'd4,	5'd5};
	rom[ 1244 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1245 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1246 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1247 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1248 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1249 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1250 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1251 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1252 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1253 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1254 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1255 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1256 ] = { 5'd3,	5'd13,	5'd2,	5'd9};
	rom[ 1257 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1258 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1259 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1260 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1261 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1262 ] = { 5'd10,	5'd12,	5'd10,	5'd2};
	rom[ 1263 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1264 ] = { 5'd9,	5'd11,	5'd3,	5'd6};
	rom[ 1265 ] = { 5'd6,	5'd11,	5'd9,	5'd11};
	rom[ 1266 ] = { 5'd9,	5'd11,	5'd9,	5'd11};
	rom[ 1267 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1268 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1269 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1270 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1271 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1272 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1273 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1274 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1275 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1276 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1277 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1278 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1279 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1280 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1281 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1282 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1283 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1284 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1285 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1286 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1287 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1288 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1289 ] = { 5'd9,	5'd13,	5'd4,	5'd5};
	rom[ 1290 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1291 ] = { 5'd9,	5'd13,	5'd4,	5'd5};
	rom[ 1292 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1293 ] = { 5'd9,	5'd13,	5'd4,	5'd5};
	rom[ 1294 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1295 ] = { 5'd10,	5'd15,	5'd2,	5'd9};
	rom[ 1296 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1297 ] = { 5'd9,	5'd13,	5'd4,	5'd5};
	rom[ 1298 ] = { 5'd11,	5'd13,	5'd4,	5'd5};
	rom[ 1299 ] = { 5'd11,	5'd17,	5'd3,	5'd7};
	rom[ 1300 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1301 ] = { 5'd6,	5'd15,	5'd6,	5'd3};
	rom[ 1302 ] = { 5'd10,	5'd12,	5'd9,	5'd3};
	rom[ 1303 ] = { 5'd16,	5'd19,	5'd4,	5'd5};
	rom[ 1304 ] = { 5'd11,	5'd13,	5'd11,	5'd4};
	rom[ 1305 ] = { 5'd8,	5'd21,	5'd6,	5'd3};
	rom[ 1306 ] = { 5'd10,	5'd15,	5'd10,	5'd9};
	rom[ 1307 ] = { 5'd3,	5'd12,	5'd10,	5'd6};
	rom[ 1308 ] = { 5'd5,	5'd20,	5'd5,	5'd4};
	rom[ 1309 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1310 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1311 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1312 ] = { 5'd12,	5'd9,	5'd11,	5'd2};
	rom[ 1313 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1314 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1315 ] = { 5'd12,	5'd14,	5'd5,	5'd4};
	rom[ 1316 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1317 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1318 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1319 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1320 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1321 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1322 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1323 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1324 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1325 ] = { 5'd15,	5'd6,	5'd4,	5'd6};
	rom[ 1326 ] = { 5'd4,	5'd6,	5'd4,	5'd6};
	rom[ 1327 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1328 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1329 ] = { 5'd14,	5'd14,	5'd3,	5'd6};
	rom[ 1330 ] = { 5'd7,	5'd14,	5'd3,	5'd6};
	rom[ 1331 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1332 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1333 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1334 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1335 ] = { 5'd11,	5'd19,	5'd6,	5'd4};
	rom[ 1336 ] = { 5'd12,	5'd4,	5'd12,	5'd2};
	rom[ 1337 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1338 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1339 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1340 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1341 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1342 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1343 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1344 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1345 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1346 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1347 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1348 ] = { 5'd12,	5'd18,	5'd3,	5'd6};
	rom[ 1349 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1350 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1351 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1352 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1353 ] = { 5'd4,	5'd16,	5'd9,	5'd2};
	rom[ 1354 ] = { 5'd10,	5'd14,	5'd3,	5'd7};
	rom[ 1355 ] = { 5'd7,	5'd16,	5'd6,	5'd3};
	rom[ 1356 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1357 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1358 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1359 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1360 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1361 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1362 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1363 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1364 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1365 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1366 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1367 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1368 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1369 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1370 ] = { 5'd7,	5'd19,	5'd6,	5'd4};
	rom[ 1371 ] = { 5'd15,	5'd17,	5'd4,	5'd7};
	rom[ 1372 ] = { 5'd5,	5'd16,	5'd4,	5'd7};
	rom[ 1373 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1374 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1375 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1376 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1377 ] = { 5'd10,	5'd9,	5'd4,	5'd5};
	rom[ 1378 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1379 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1380 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1381 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1382 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1383 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1384 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1385 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1386 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1387 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1388 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1389 ] = { 5'd9,	5'd7,	5'd5,	5'd4};
	rom[ 1390 ] = { 5'd10,	5'd7,	5'd5,	5'd4};
	rom[ 1391 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1392 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1393 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1394 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1395 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1396 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1397 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1398 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1399 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1400 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1401 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1402 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1403 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1404 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1405 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1406 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1407 ] = { 5'd10,	5'd12,	5'd4,	5'd5};
	rom[ 1408 ] = { 5'd14,	5'd7,	5'd3,	5'd7};
	rom[ 1409 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1410 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1411 ] = { 5'd12,	5'd11,	5'd6,	5'd4};
	rom[ 1412 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1413 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1414 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1415 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1416 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1417 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1418 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1419 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1420 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1421 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1422 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1423 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1424 ] = { 5'd7,	5'd15,	5'd5,	5'd4};
	rom[ 1425 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1426 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1427 ] = { 5'd10,	5'd13,	5'd8,	5'd4};
	rom[ 1428 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1429 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1430 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1431 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1432 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1433 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1434 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1435 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1436 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1437 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1438 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1439 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1440 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1441 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1442 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1443 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1444 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1445 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1446 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1447 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1448 ] = { 5'd1,	5'd18,	5'd11,	5'd2};
	rom[ 1449 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1450 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1451 ] = { 5'd8,	5'd21,	5'd6,	5'd3};
	rom[ 1452 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1453 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1454 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1455 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1456 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1457 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1458 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1459 ] = { 5'd7,	5'd21,	5'd6,	5'd3};
	rom[ 1460 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1461 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1462 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1463 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1464 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1465 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1466 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1467 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1468 ] = { 5'd17,	5'd7,	5'd3,	5'd7};
	rom[ 1469 ] = { 5'd4,	5'd7,	5'd3,	5'd7};
	rom[ 1470 ] = { 5'd14,	5'd8,	5'd3,	5'd8};
	rom[ 1471 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1472 ] = { 5'd3,	5'd20,	5'd9,	5'd3};
	rom[ 1473 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1474 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1475 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1476 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1477 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1478 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1479 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1480 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1481 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1482 ] = { 5'd6,	5'd6,	5'd6,	5'd6};
	rom[ 1483 ] = { 5'd12,	5'd16,	5'd4,	5'd6};
	rom[ 1484 ] = { 5'd14,	5'd20,	5'd5,	5'd4};
	rom[ 1485 ] = { 5'd5,	5'd20,	5'd5,	5'd4};
	rom[ 1486 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1487 ] = { 5'd11,	5'd20,	5'd5,	5'd4};
	rom[ 1488 ] = { 5'd7,	5'd9,	5'd6,	5'd3};
	rom[ 1489 ] = { 5'd11,	5'd15,	5'd2,	5'd9};
	rom[ 1490 ] = { 5'd10,	5'd16,	5'd3,	5'd7};
	rom[ 1491 ] = { 5'd11,	5'd16,	5'd3,	5'd7};
	rom[ 1492 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1493 ] = { 5'd7,	5'd16,	5'd3,	5'd8};
	rom[ 1494 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1495 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1496 ] = { 5'd10,	5'd10,	5'd4,	5'd9};
	rom[ 1497 ] = { 5'd10,	5'd9,	5'd8,	5'd4};
	rom[ 1498 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1499 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1500 ] = { 5'd15,	5'd14,	5'd4,	5'd10};
	rom[ 1501 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1502 ] = { 5'd15,	5'd14,	5'd4,	5'd10};
	rom[ 1503 ] = { 5'd5,	5'd14,	5'd4,	5'd10};
	rom[ 1504 ] = { 5'd11,	5'd15,	5'd4,	5'd7};
	rom[ 1505 ] = { 5'd9,	5'd15,	5'd4,	5'd7};
	rom[ 1506 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1507 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1508 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1509 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1510 ] = { 5'd10,	5'd10,	5'd4,	5'd8};
	rom[ 1511 ] = { 5'd12,	5'd5,	5'd12,	5'd3};
	rom[ 1512 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1513 ] = { 5'd7,	5'd8,	5'd6,	5'd6};
	rom[ 1514 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1515 ] = { 5'd8,	5'd8,	5'd4,	5'd5};
	rom[ 1516 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1517 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1518 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1519 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1520 ] = { 5'd12,	5'd11,	5'd6,	5'd3};
	rom[ 1521 ] = { 5'd6,	5'd11,	5'd6,	5'd3};
	rom[ 1522 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1523 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1524 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1525 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1526 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1527 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1528 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1529 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1530 ] = { 5'd9,	5'd16,	5'd6,	5'd5};
	rom[ 1531 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1532 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1533 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1534 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1535 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1536 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1537 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1538 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1539 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1540 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1541 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1542 ] = { 5'd4,	5'd11,	5'd8,	5'd6};
	rom[ 1543 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1544 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1545 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1546 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1547 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1548 ] = { 5'd16,	5'd7,	5'd3,	5'd6};
	rom[ 1549 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1550 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1551 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1552 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1553 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1554 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1555 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1556 ] = { 5'd10,	5'd10,	5'd4,	5'd5};
	rom[ 1557 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1558 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1559 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1560 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1561 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1562 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1563 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1564 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1565 ] = { 5'd9,	5'd21,	5'd6,	5'd3};
	rom[ 1566 ] = { 5'd12,	5'd11,	5'd10,	5'd3};
	rom[ 1567 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1568 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1569 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1570 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1571 ] = { 5'd0,	5'd4,	5'd12,	5'd3};
	rom[ 1572 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1573 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1574 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1575 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1576 ] = { 5'd12,	5'd9,	5'd7,	5'd3};
	rom[ 1577 ] = { 5'd13,	5'd10,	5'd4,	5'd5};
	rom[ 1578 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1579 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1580 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1581 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1582 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1583 ] = { 5'd8,	5'd8,	5'd4,	5'd5};
	rom[ 1584 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1585 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1586 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1587 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1588 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1589 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1590 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1591 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1592 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1593 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1594 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1595 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1596 ] = { 5'd6,	5'd11,	5'd6,	5'd3};
	rom[ 1597 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1598 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1599 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1600 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1601 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1602 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1603 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1604 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1605 ] = { 5'd9,	5'd21,	5'd6,	5'd3};
	rom[ 1606 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1607 ] = { 5'd16,	5'd18,	5'd4,	5'd5};
	rom[ 1608 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1609 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1610 ] = { 5'd4,	5'd18,	5'd4,	5'd5};
	rom[ 1611 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1612 ] = { 5'd11,	5'd6,	5'd6,	5'd4};
	rom[ 1613 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1614 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1615 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1616 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1617 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1618 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1619 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1620 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1621 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1622 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1623 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1624 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1625 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1626 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1627 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1628 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1629 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1630 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1631 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1632 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1633 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1634 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1635 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1636 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1637 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1638 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1639 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1640 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1641 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1642 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1643 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1644 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1645 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1646 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1647 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1648 ] = { 5'd10,	5'd10,	5'd5,	5'd4};
	rom[ 1649 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1650 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1651 ] = { 5'd2,	5'd12,	5'd11,	5'd7};
	rom[ 1652 ] = { 5'd7,	5'd15,	5'd4,	5'd5};
	rom[ 1653 ] = { 5'd17,	5'd6,	5'd3,	5'd6};
	rom[ 1654 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1655 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1656 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1657 ] = { 5'd15,	5'd18,	5'd4,	5'd5};
	rom[ 1658 ] = { 5'd4,	5'd6,	5'd3,	5'd6};
	rom[ 1659 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1660 ] = { 5'd5,	5'd18,	5'd4,	5'd5};
	rom[ 1661 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1662 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1663 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1664 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1665 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1666 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1667 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1668 ] = { 5'd10,	5'd5,	5'd5,	5'd4};
	rom[ 1669 ] = { 5'd11,	5'd21,	5'd6,	5'd3};
	rom[ 1670 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1671 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1672 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1673 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1674 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1675 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1676 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1677 ] = { 5'd6,	5'd7,	5'd9,	5'd3};
	rom[ 1678 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1679 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1680 ] = { 5'd11,	5'd12,	5'd11,	5'd8};
	rom[ 1681 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1682 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1683 ] = { 5'd12,	5'd9,	5'd6,	5'd9};
	rom[ 1684 ] = { 5'd6,	5'd9,	5'd6,	5'd9};
	rom[ 1685 ] = { 5'd1,	5'd3,	5'd11,	5'd2};
	rom[ 1686 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1687 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1688 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1689 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1690 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1691 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1692 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1693 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1694 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1695 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1696 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1697 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1698 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1699 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1700 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1701 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1702 ] = { 5'd10,	5'd10,	5'd5,	5'd4};
	rom[ 1703 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1704 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1705 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1706 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1707 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1708 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1709 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1710 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1711 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1712 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1713 ] = { 5'd0,	5'd12,	5'd12,	5'd3};
	rom[ 1714 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1715 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1716 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1717 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1718 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1719 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1720 ] = { 5'd7,	5'd21,	5'd6,	5'd3};
	rom[ 1721 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1722 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1723 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1724 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1725 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1726 ] = { 5'd12,	5'd12,	5'd5,	5'd5};
	rom[ 1727 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1728 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1729 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1730 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1731 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1732 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1733 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1734 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1735 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1736 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1737 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1738 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1739 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1740 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1741 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1742 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1743 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1744 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1745 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1746 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1747 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1748 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1749 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1750 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1751 ] = { 5'd11,	5'd16,	5'd7,	5'd6};
	rom[ 1752 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1753 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1754 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1755 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1756 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1757 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1758 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1759 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1760 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1761 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1762 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1763 ] = { 5'd12,	5'd8,	5'd8,	5'd8};
	rom[ 1764 ] = { 5'd6,	5'd9,	5'd7,	5'd3};
	rom[ 1765 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1766 ] = { 5'd9,	5'd19,	5'd6,	5'd4};
	rom[ 1767 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1768 ] = { 5'd5,	5'd9,	5'd7,	5'd3};
	rom[ 1769 ] = { 5'd12,	5'd11,	5'd9,	5'd5};
	rom[ 1770 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1771 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1772 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1773 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1774 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1775 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1776 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1777 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1778 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1779 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1780 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1781 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1782 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1783 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1784 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1785 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1786 ] = { 5'd14,	5'd16,	5'd3,	5'd7};
	rom[ 1787 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1788 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1789 ] = { 5'd7,	5'd9,	5'd6,	5'd5};
	rom[ 1790 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1791 ] = { 5'd5,	5'd7,	5'd4,	5'd5};
	rom[ 1792 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1793 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1794 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1795 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1796 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1797 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1798 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1799 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1800 ] = { 5'd10,	5'd15,	5'd2,	5'd9};
	rom[ 1801 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1802 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1803 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1804 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1805 ] = { 5'd11,	5'd7,	5'd4,	5'd5};
	rom[ 1806 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1807 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1808 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1809 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1810 ] = { 5'd5,	5'd9,	5'd8,	5'd3};
	rom[ 1811 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1812 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1813 ] = { 5'd12,	5'd11,	5'd12,	5'd11};
	rom[ 1814 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1815 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1816 ] = { 5'd1,	5'd21,	5'd11,	5'd2};
	rom[ 1817 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1818 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1819 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1820 ] = { 5'd10,	5'd21,	5'd6,	5'd3};
	rom[ 1821 ] = { 5'd8,	5'd21,	5'd6,	5'd3};
	rom[ 1822 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1823 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1824 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1825 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1826 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1827 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1828 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1829 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1830 ] = { 5'd0,	5'd7,	5'd12,	5'd2};
	rom[ 1831 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1832 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1833 ] = { 5'd3,	5'd18,	5'd3,	5'd6};
	rom[ 1834 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1835 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1836 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1837 ] = { 5'd12,	5'd10,	5'd5,	5'd4};
	rom[ 1838 ] = { 5'd6,	5'd9,	5'd7,	5'd3};
	rom[ 1839 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1840 ] = { 5'd14,	5'd16,	5'd3,	5'd6};
	rom[ 1841 ] = { 5'd7,	5'd16,	5'd3,	5'd6};
	rom[ 1842 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1843 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1844 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1845 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1846 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1847 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1848 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1849 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1850 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1851 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1852 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1853 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1854 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1855 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1856 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1857 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1858 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1859 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1860 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1861 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1862 ] = { 5'd8,	5'd15,	5'd4,	5'd5};
	rom[ 1863 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1864 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1865 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1866 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1867 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1868 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1869 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1870 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1871 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1872 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1873 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1874 ] = { 5'd8,	5'd5,	5'd6,	5'd3};
	rom[ 1875 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1876 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1877 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1878 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1879 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1880 ] = { 5'd14,	5'd9,	5'd3,	5'd6};
	rom[ 1881 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1882 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1883 ] = { 5'd7,	5'd9,	5'd3,	5'd6};
	rom[ 1884 ] = { 5'd12,	5'd11,	5'd6,	5'd3};
	rom[ 1885 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1886 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1887 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1888 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1889 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1890 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1891 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1892 ] = { 5'd9,	5'd9,	5'd5,	5'd4};
	rom[ 1893 ] = { 5'd12,	5'd8,	5'd8,	5'd4};
	rom[ 1894 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1895 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1896 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1897 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1898 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1899 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1900 ] = { 5'd10,	5'd16,	5'd7,	5'd3};
	rom[ 1901 ] = { 5'd7,	5'd16,	5'd7,	5'd3};
	rom[ 1902 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1903 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1904 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1905 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1906 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1907 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1908 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1909 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1910 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1911 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1912 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1913 ] = { 5'd9,	5'd10,	5'd9,	5'd2};
	rom[ 1914 ] = { 5'd3,	5'd13,	5'd10,	5'd3};
	rom[ 1915 ] = { 5'd11,	5'd13,	5'd10,	5'd3};
	rom[ 1916 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1917 ] = { 5'd11,	5'd16,	5'd10,	5'd4};
	rom[ 1918 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1919 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1920 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1921 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1922 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1923 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1924 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1925 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1926 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1927 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1928 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1929 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1930 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1931 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1932 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1933 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1934 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1935 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1936 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1937 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1938 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1939 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1940 ] = { 5'd11,	5'd14,	5'd3,	5'd7};
	rom[ 1941 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1942 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1943 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1944 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1945 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1946 ] = { 5'd6,	5'd9,	5'd6,	5'd3};
	rom[ 1947 ] = { 5'd12,	5'd21,	5'd10,	5'd2};
	rom[ 1948 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1949 ] = { 5'd12,	5'd12,	5'd9,	5'd7};
	rom[ 1950 ] = { 5'd15,	5'd15,	5'd2,	5'd9};
	rom[ 1951 ] = { 5'd7,	5'd15,	5'd2,	5'd9};
	rom[ 1952 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1953 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1954 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1955 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1956 ] = { 5'd4,	5'd4,	5'd8,	5'd3};
	rom[ 1957 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1958 ] = { 5'd17,	5'd7,	5'd3,	5'd6};
	rom[ 1959 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1960 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1961 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1962 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1963 ] = { 5'd4,	5'd7,	5'd3,	5'd6};
	rom[ 1964 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1965 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1966 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1967 ] = { 5'd7,	5'd8,	5'd6,	5'd3};
	rom[ 1968 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1969 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1970 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1971 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1972 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1973 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1974 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1975 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1976 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1977 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1978 ] = { 5'd5,	5'd12,	5'd9,	5'd3};
	rom[ 1979 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1980 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1981 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1982 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1983 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1984 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1985 ] = { 5'd7,	5'd21,	5'd6,	5'd3};
	rom[ 1986 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1987 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1988 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1989 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1990 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1991 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1992 ] = { 5'd4,	5'd12,	5'd10,	5'd3};
	rom[ 1993 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1994 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1995 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1996 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1997 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1998 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 1999 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2000 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2001 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2002 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2003 ] = { 5'd11,	5'd9,	5'd8,	5'd3};
	rom[ 2004 ] = { 5'd5,	5'd11,	5'd8,	5'd7};
	rom[ 2005 ] = { 5'd12,	5'd2,	5'd12,	5'd2};
	rom[ 2006 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2007 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2008 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2009 ] = { 5'd12,	5'd8,	5'd4,	5'd5};
	rom[ 2010 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2011 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2012 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2013 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2014 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2015 ] = { 5'd12,	5'd18,	5'd12,	5'd2};
	rom[ 2016 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2017 ] = { 5'd5,	5'd17,	5'd4,	5'd7};
	rom[ 2018 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2019 ] = { 5'd11,	5'd12,	5'd5,	5'd12};
	rom[ 2020 ] = { 5'd7,	5'd12,	5'd7,	5'd7};
	rom[ 2021 ] = { 5'd12,	5'd12,	5'd5,	5'd4};
	rom[ 2022 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2023 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2024 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2025 ] = { 5'd12,	5'd15,	5'd11,	5'd2};
	rom[ 2026 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2027 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2028 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2029 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2030 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2031 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2032 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2033 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2034 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2035 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2036 ] = { 5'd13,	5'd12,	5'd2,	5'd11};
	rom[ 2037 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2038 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2039 ] = { 5'd12,	5'd14,	5'd9,	5'd2};
	rom[ 2040 ] = { 5'd13,	5'd12,	5'd2,	5'd11};
	rom[ 2041 ] = { 5'd9,	5'd12,	5'd2,	5'd11};
	rom[ 2042 ] = { 5'd4,	5'd9,	5'd10,	5'd2};
	rom[ 2043 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2044 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2045 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2046 ] = { 5'd15,	5'd6,	5'd4,	5'd6};
	rom[ 2047 ] = { 5'd5,	5'd6,	5'd4,	5'd6};
	rom[ 2048 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2049 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2050 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2051 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2052 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2053 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2054 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2055 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2056 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2057 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2058 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2059 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2060 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2061 ] = { 5'd3,	5'd17,	5'd3,	5'd7};
	rom[ 2062 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2063 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2064 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2065 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2066 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2067 ] = { 5'd9,	5'd11,	5'd5,	5'd5};
	rom[ 2068 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2069 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2070 ] = { 5'd11,	5'd11,	5'd2,	5'd10};
	rom[ 2071 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2072 ] = { 5'd11,	5'd11,	5'd2,	5'd10};
	rom[ 2073 ] = { 5'd6,	5'd20,	5'd5,	5'd4};
	rom[ 2074 ] = { 5'd11,	5'd11,	5'd2,	5'd10};
	rom[ 2075 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2076 ] = { 5'd11,	5'd11,	5'd2,	5'd10};
	rom[ 2077 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2078 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2079 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2080 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2081 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2082 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2083 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2084 ] = { 5'd6,	5'd2,	5'd9,	5'd2};
	rom[ 2085 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2086 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2087 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2088 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2089 ] = { 5'd12,	5'd15,	5'd2,	5'd9};
	rom[ 2090 ] = { 5'd11,	5'd11,	5'd2,	5'd10};
	rom[ 2091 ] = { 5'd11,	5'd11,	5'd2,	5'd10};
	rom[ 2092 ] = { 5'd5,	5'd12,	5'd9,	5'd3};
	rom[ 2093 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2094 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2095 ] = { 5'd9,	5'd4,	5'd9,	5'd4};
	rom[ 2096 ] = { 5'd6,	5'd11,	5'd7,	5'd6};
	rom[ 2097 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2098 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2099 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2100 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2101 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2102 ] = { 5'd13,	5'd8,	5'd3,	5'd6};
	rom[ 2103 ] = { 5'd12,	5'd15,	5'd2,	5'd9};
	rom[ 2104 ] = { 5'd7,	5'd16,	5'd5,	5'd8};
	rom[ 2105 ] = { 5'd12,	5'd7,	5'd4,	5'd6};
	rom[ 2106 ] = { 5'd7,	5'd8,	5'd6,	5'd7};
	rom[ 2107 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2108 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2109 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2110 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2111 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2112 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2113 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2114 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2115 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2116 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2117 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2118 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2119 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2120 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2121 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2122 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2123 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2124 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2125 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2126 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2127 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2128 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2129 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2130 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2131 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2132 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2133 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2134 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2135 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2136 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2137 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2138 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2139 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2140 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2141 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2142 ] = { 5'd11,	5'd13,	5'd6,	5'd7};
	rom[ 2143 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2144 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2145 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2146 ] = { 5'd10,	5'd11,	5'd6,	5'd10};
	rom[ 2147 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2148 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2149 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2150 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2151 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2152 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2153 ] = { 5'd19,	5'd13,	5'd2,	5'd9};
	rom[ 2154 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2155 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2156 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2157 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2158 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2159 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2160 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2161 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2162 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2163 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2164 ] = { 5'd12,	5'd18,	5'd3,	5'd6};
	rom[ 2165 ] = { 5'd14,	5'd19,	5'd4,	5'd5};
	rom[ 2166 ] = { 5'd6,	5'd19,	5'd4,	5'd5};
	rom[ 2167 ] = { 5'd10,	5'd21,	5'd6,	5'd3};
	rom[ 2168 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2169 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2170 ] = { 5'd11,	5'd9,	5'd7,	5'd3};
	rom[ 2171 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2172 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2173 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2174 ] = { 5'd10,	5'd15,	5'd3,	5'd7};
	rom[ 2175 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2176 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2177 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2178 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2179 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2180 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2181 ] = { 5'd16,	5'd5,	5'd4,	5'd5};
	rom[ 2182 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2183 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2184 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2185 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2186 ] = { 5'd4,	5'd5,	5'd4,	5'd5};
	rom[ 2187 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2188 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2189 ] = { 5'd3,	5'd5,	5'd9,	5'd5};
	rom[ 2190 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2191 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2192 ] = { 5'd6,	5'd12,	5'd6,	5'd3};
	rom[ 2193 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2194 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2195 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2196 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2197 ] = { 5'd19,	5'd13,	5'd2,	5'd9};
	rom[ 2198 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2199 ] = { 5'd19,	5'd13,	5'd2,	5'd9};
	rom[ 2200 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2201 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2202 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2203 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2204 ] = { 5'd3,	5'd14,	5'd2,	5'd9};
	rom[ 2205 ] = { 5'd9,	5'd13,	5'd4,	5'd5};
	rom[ 2206 ] = { 5'd11,	5'd13,	5'd4,	5'd5};
	rom[ 2207 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2208 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2209 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2210 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2211 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2212 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2213 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2214 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2215 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2216 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2217 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2218 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2219 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2220 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2221 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2222 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2223 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2224 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2225 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2226 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2227 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2228 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2229 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2230 ] = { 5'd5,	5'd14,	5'd2,	5'd10};
	rom[ 2231 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2232 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2233 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2234 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2235 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2236 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2237 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2238 ] = { 5'd6,	5'd10,	5'd3,	5'd6};
	rom[ 2239 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2240 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2241 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2242 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2243 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2244 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2245 ] = { 5'd13,	5'd15,	5'd4,	5'd5};
	rom[ 2246 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2247 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2248 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2249 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2250 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2251 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2252 ] = { 5'd7,	5'd15,	5'd4,	5'd5};
	rom[ 2253 ] = { 5'd8,	5'd21,	5'd8,	5'd3};
	rom[ 2254 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2255 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2256 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2257 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2258 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2259 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2260 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2261 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2262 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2263 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2264 ] = { 5'd12,	5'd17,	5'd3,	5'd6};
	rom[ 2265 ] = { 5'd0,	5'd9,	5'd12,	5'd4};
	rom[ 2266 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2267 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2268 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2269 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2270 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2271 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2272 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2273 ] = { 5'd6,	5'd13,	5'd6,	5'd4};
	rom[ 2274 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2275 ] = { 5'd11,	5'd10,	5'd6,	5'd8};
	rom[ 2276 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2277 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2278 ] = { 5'd11,	5'd14,	5'd11,	5'd2};
	rom[ 2279 ] = { 5'd1,	5'd15,	5'd11,	5'd3};
	rom[ 2280 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2281 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2282 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2283 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2284 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2285 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2286 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2287 ] = { 5'd10,	5'd20,	5'd5,	5'd4};
	rom[ 2288 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2289 ] = { 5'd12,	5'd16,	5'd3,	5'd6};
	rom[ 2290 ] = { 5'd9,	5'd16,	5'd3,	5'd6};
	rom[ 2291 ] = { 5'd16,	5'd18,	5'd3,	5'd6};
	rom[ 2292 ] = { 5'd5,	5'd18,	5'd3,	5'd6};
	rom[ 2293 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2294 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2295 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2296 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2297 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2298 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2299 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2300 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2301 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2302 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2303 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2304 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2305 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2306 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2307 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2308 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2309 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2310 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2311 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2312 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2313 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2314 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2315 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2316 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2317 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2318 ] = { 5'd13,	5'd14,	5'd4,	5'd5};
	rom[ 2319 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2320 ] = { 5'd13,	5'd14,	5'd4,	5'd5};
	rom[ 2321 ] = { 5'd12,	5'd16,	5'd5,	5'd5};
	rom[ 2322 ] = { 5'd4,	5'd15,	5'd9,	5'd2};
	rom[ 2323 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2324 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2325 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2326 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2327 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2328 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2329 ] = { 5'd9,	5'd21,	5'd6,	5'd3};
	rom[ 2330 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2331 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2332 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2333 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2334 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2335 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2336 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2337 ] = { 5'd8,	5'd15,	5'd2,	5'd9};
	rom[ 2338 ] = { 5'd14,	5'd15,	5'd3,	5'd6};
	rom[ 2339 ] = { 5'd7,	5'd15,	5'd3,	5'd6};
	rom[ 2340 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2341 ] = { 5'd9,	5'd22,	5'd9,	5'd2};
	rom[ 2342 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2343 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2344 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2345 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2346 ] = { 5'd19,	5'd13,	5'd2,	5'd11};
	rom[ 2347 ] = { 5'd3,	5'd13,	5'd2,	5'd11};
	rom[ 2348 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2349 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2350 ] = { 5'd11,	5'd15,	5'd2,	5'd9};
	rom[ 2351 ] = { 5'd12,	5'd16,	5'd5,	5'd7};
	rom[ 2352 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2353 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2354 ] = { 5'd20,	5'd14,	5'd2,	5'd10};
	rom[ 2355 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2356 ] = { 5'd7,	5'd7,	5'd5,	5'd7};
	rom[ 2357 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2358 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2359 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2360 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2361 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2362 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2363 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2364 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2365 ] = { 5'd8,	5'd20,	5'd5,	5'd4};
	rom[ 2366 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2367 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2368 ] = { 5'd20,	5'd14,	5'd2,	5'd10};
	rom[ 2369 ] = { 5'd2,	5'd14,	5'd2,	5'd10};
	rom[ 2370 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2371 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2372 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2373 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2374 ] = { 5'd7,	5'd12,	5'd7,	5'd10};
	rom[ 2375 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2376 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2377 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2378 ] = { 5'd7,	5'd11,	5'd8,	5'd10};
	rom[ 2379 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2380 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2381 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2382 ] = { 5'd7,	5'd11,	5'd8,	5'd10};
	rom[ 2383 ] = { 5'd9,	5'd11,	5'd8,	5'd10};
	rom[ 2384 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2385 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2386 ] = { 5'd7,	5'd10,	5'd5,	5'd4};
	rom[ 2387 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2388 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2389 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2390 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2391 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2392 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2393 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2394 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2395 ] = { 5'd12,	5'd15,	5'd2,	5'd9};
	rom[ 2396 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2397 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2398 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2399 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2400 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2401 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2402 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2403 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2404 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2405 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2406 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2407 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2408 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2409 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2410 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2411 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2412 ] = { 5'd2,	5'd4,	5'd10,	5'd2};
	rom[ 2413 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2414 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2415 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2416 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2417 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2418 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2419 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2420 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2421 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2422 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2423 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2424 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2425 ] = { 5'd12,	5'd14,	5'd10,	5'd2};
	rom[ 2426 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2427 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2428 ] = { 5'd15,	5'd12,	5'd2,	5'd11};
	rom[ 2429 ] = { 5'd7,	5'd12,	5'd2,	5'd11};
	rom[ 2430 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2431 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2432 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2433 ] = { 5'd11,	5'd11,	5'd6,	5'd3};
	rom[ 2434 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2435 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2436 ] = { 5'd12,	5'd12,	5'd3,	5'd6};
	rom[ 2437 ] = { 5'd9,	5'd12,	5'd3,	5'd6};
	rom[ 2438 ] = { 5'd5,	5'd13,	5'd7,	5'd4};
	rom[ 2439 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2440 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2441 ] = { 5'd6,	5'd14,	5'd2,	5'd9};
	rom[ 2442 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2443 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2444 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2445 ] = { 5'd12,	5'd17,	5'd3,	5'd7};
	rom[ 2446 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2447 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2448 ] = { 5'd1,	5'd11,	5'd11,	5'd7};
	rom[ 2449 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2450 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2451 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2452 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2453 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2454 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2455 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2456 ] = { 5'd4,	5'd15,	5'd9,	5'd2};
	rom[ 2457 ] = { 5'd11,	5'd15,	5'd9,	5'd2};
	rom[ 2458 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2459 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2460 ] = { 5'd6,	5'd12,	5'd9,	5'd12};
	rom[ 2461 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2462 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2463 ] = { 5'd10,	5'd12,	5'd9,	5'd3};
	rom[ 2464 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2465 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2466 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2467 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2468 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2469 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2470 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2471 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2472 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2473 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2474 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2475 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2476 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2477 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2478 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2479 ] = { 5'd12,	5'd12,	5'd6,	5'd7};
	rom[ 2480 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2481 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2482 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2483 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2484 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2485 ] = { 5'd12,	5'd11,	5'd4,	5'd5};
	rom[ 2486 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2487 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2488 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2489 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2490 ] = { 5'd13,	5'd19,	5'd5,	5'd4};
	rom[ 2491 ] = { 5'd3,	5'd7,	5'd3,	5'd6};
	rom[ 2492 ] = { 5'd10,	5'd6,	5'd3,	5'd6};
	rom[ 2493 ] = { 5'd12,	5'd6,	5'd5,	5'd6};
	rom[ 2494 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2495 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2496 ] = { 5'd6,	5'd11,	5'd9,	5'd2};
	rom[ 2497 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2498 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2499 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2500 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2501 ] = { 5'd7,	5'd10,	5'd4,	5'd10};
	rom[ 2502 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2503 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2504 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2505 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2506 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2507 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2508 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2509 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2510 ] = { 5'd12,	5'd3,	5'd6,	5'd3};
	rom[ 2511 ] = { 5'd4,	5'd9,	5'd9,	5'd2};
	rom[ 2512 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2513 ] = { 5'd7,	5'd15,	5'd5,	5'd6};
	rom[ 2514 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2515 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2516 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2517 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2518 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2519 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2520 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2521 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2522 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2523 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2524 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2525 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2526 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2527 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2528 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2529 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2530 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2531 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2532 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2533 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2534 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2535 ] = { 5'd18,	5'd11,	5'd3,	5'd10};
	rom[ 2536 ] = { 5'd3,	5'd11,	5'd3,	5'd10};
	rom[ 2537 ] = { 5'd13,	5'd12,	5'd2,	5'd9};
	rom[ 2538 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2539 ] = { 5'd12,	5'd12,	5'd6,	5'd3};
	rom[ 2540 ] = { 5'd9,	5'd12,	5'd2,	5'd9};
	rom[ 2541 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2542 ] = { 5'd6,	5'd12,	5'd6,	5'd3};
	rom[ 2543 ] = { 5'd14,	5'd14,	5'd4,	5'd10};
	rom[ 2544 ] = { 5'd6,	5'd14,	5'd4,	5'd10};
	rom[ 2545 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2546 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2547 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2548 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2549 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2550 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2551 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2552 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2553 ] = { 5'd5,	5'd9,	5'd7,	5'd3};
	rom[ 2554 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2555 ] = { 5'd6,	5'd14,	5'd6,	5'd3};
	rom[ 2556 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2557 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2558 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2559 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2560 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2561 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2562 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2563 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2564 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2565 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2566 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2567 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2568 ] = { 5'd9,	5'd10,	5'd9,	5'd7};
	rom[ 2569 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2570 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2571 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2572 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2573 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2574 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2575 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2576 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2577 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2578 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2579 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2580 ] = { 5'd12,	5'd15,	5'd3,	5'd9};
	rom[ 2581 ] = { 5'd15,	5'd19,	5'd4,	5'd5};
	rom[ 2582 ] = { 5'd5,	5'd19,	5'd4,	5'd5};
	rom[ 2583 ] = { 5'd11,	5'd5,	5'd4,	5'd5};
	rom[ 2584 ] = { 5'd9,	5'd5,	5'd4,	5'd5};
	rom[ 2585 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2586 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2587 ] = { 5'd2,	5'd11,	5'd10,	5'd3};
	rom[ 2588 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2589 ] = { 5'd10,	5'd13,	5'd4,	5'd8};
	rom[ 2590 ] = { 5'd11,	5'd13,	5'd8,	5'd4};
	rom[ 2591 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2592 ] = { 5'd12,	5'd16,	5'd5,	5'd4};
	rom[ 2593 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2594 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2595 ] = { 5'd13,	5'd8,	5'd5,	5'd4};
	rom[ 2596 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2597 ] = { 5'd8,	5'd13,	5'd5,	5'd6};
	rom[ 2598 ] = { 5'd11,	5'd13,	5'd5,	5'd6};
	rom[ 2599 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2600 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2601 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2602 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2603 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2604 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2605 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2606 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2607 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2608 ] = { 5'd12,	5'd12,	5'd9,	5'd3};
	rom[ 2609 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2610 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2611 ] = { 5'd4,	5'd9,	5'd9,	5'd2};
	rom[ 2612 ] = { 5'd8,	5'd11,	5'd6,	5'd10};
	rom[ 2613 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2614 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2615 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2616 ] = { 5'd10,	5'd9,	5'd10,	5'd3};
	rom[ 2617 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2618 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2619 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2620 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2621 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2622 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2623 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2624 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2625 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2626 ] = { 5'd8,	5'd19,	5'd4,	5'd5};
	rom[ 2627 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2628 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2629 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2630 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2631 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2632 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2633 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2634 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2635 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2636 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2637 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2638 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2639 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2640 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2641 ] = { 5'd9,	5'd13,	5'd5,	5'd7};
	rom[ 2642 ] = { 5'd5,	5'd11,	5'd4,	5'd5};
	rom[ 2643 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2644 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2645 ] = { 5'd7,	5'd15,	5'd7,	5'd7};
	rom[ 2646 ] = { 5'd10,	5'd15,	5'd7,	5'd7};
	rom[ 2647 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2648 ] = { 5'd6,	5'd8,	5'd3,	5'd6};
	rom[ 2649 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2650 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2651 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2652 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2653 ] = { 5'd0,	5'd14,	5'd12,	5'd5};
	rom[ 2654 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2655 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2656 ] = { 5'd9,	5'd3,	5'd9,	5'd2};
	rom[ 2657 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2658 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2659 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2660 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2661 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2662 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2663 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2664 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2665 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2666 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2667 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2668 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2669 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2670 ] = { 5'd12,	5'd13,	5'd8,	5'd10};
	rom[ 2671 ] = { 5'd7,	5'd12,	5'd5,	5'd6};
	rom[ 2672 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2673 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2674 ] = { 5'd10,	5'd11,	5'd6,	5'd4};
	rom[ 2675 ] = { 5'd8,	5'd16,	5'd4,	5'd5};
	rom[ 2676 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2677 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2678 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2679 ] = { 5'd4,	5'd9,	5'd9,	5'd2};
	rom[ 2680 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2681 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2682 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2683 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2684 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2685 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2686 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2687 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2688 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2689 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2690 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2691 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2692 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2693 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2694 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2695 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2696 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2697 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2698 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2699 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2700 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2701 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2702 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2703 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2704 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2705 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2706 ] = { 5'd12,	5'd7,	5'd9,	5'd3};
	rom[ 2707 ] = { 5'd5,	5'd9,	5'd8,	5'd4};
	rom[ 2708 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2709 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2710 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2711 ] = { 5'd14,	5'd5,	5'd5,	5'd4};
	rom[ 2712 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2713 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2714 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2715 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2716 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2717 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2718 ] = { 5'd9,	5'd21,	5'd6,	5'd3};
	rom[ 2719 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2720 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2721 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2722 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2723 ] = { 5'd10,	5'd5,	5'd6,	5'd3};
	rom[ 2724 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2725 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2726 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2727 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2728 ] = { 5'd6,	5'd9,	5'd7,	5'd3};
	rom[ 2729 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2730 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2731 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2732 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2733 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2734 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2735 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2736 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2737 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2738 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2739 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2740 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2741 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2742 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2743 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2744 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2745 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2746 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2747 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2748 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2749 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2750 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2751 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2752 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2753 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2754 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2755 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2756 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2757 ] = { 5'd11,	5'd9,	5'd6,	5'd3};
	rom[ 2758 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2759 ] = { 5'd10,	5'd15,	5'd3,	5'd6};
	rom[ 2760 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2761 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2762 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2763 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2764 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2765 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2766 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2767 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2768 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2769 ] = { 5'd10,	5'd14,	5'd6,	5'd8};
	rom[ 2770 ] = { 5'd19,	5'd15,	5'd2,	5'd9};
	rom[ 2771 ] = { 5'd3,	5'd15,	5'd2,	5'd9};
	rom[ 2772 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2773 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2774 ] = { 5'd12,	5'd21,	5'd6,	5'd3};
	rom[ 2775 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2776 ] = { 5'd12,	5'd20,	5'd5,	5'd4};
	rom[ 2777 ] = { 5'd7,	5'd20,	5'd5,	5'd4};
	rom[ 2778 ] = { 5'd14,	5'd6,	5'd5,	5'd6};
	rom[ 2779 ] = { 5'd5,	5'd6,	5'd5,	5'd6};
	rom[ 2780 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2781 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2782 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2783 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2784 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2785 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2786 ] = { 5'd3,	5'd11,	5'd9,	5'd6};
	rom[ 2787 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2788 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2789 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2790 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2791 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2792 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2793 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2794 ] = { 5'd13,	5'd19,	5'd4,	5'd5};
	rom[ 2795 ] = { 5'd7,	5'd19,	5'd4,	5'd5};
	rom[ 2796 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2797 ] = { 5'd11,	5'd14,	5'd6,	5'd3};
	rom[ 2798 ] = { 5'd10,	5'd10,	5'd4,	5'd5};
	rom[ 2799 ] = { 5'd12,	5'd9,	5'd6,	5'd5};
	rom[ 2800 ] = { 5'd6,	5'd13,	5'd9,	5'd5};
	rom[ 2801 ] = { 5'd9,	5'd13,	5'd9,	5'd5};
	rom[ 2802 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2803 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2804 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2805 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2806 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2807 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2808 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2809 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2810 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2811 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2812 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2813 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2814 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2815 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2816 ] = { 5'd15,	5'd17,	5'd3,	5'd7};
	rom[ 2817 ] = { 5'd6,	5'd17,	5'd3,	5'd7};
	rom[ 2818 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2819 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2820 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2821 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2822 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2823 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2824 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2825 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2826 ] = { 5'd6,	5'd12,	5'd8,	5'd3};
	rom[ 2827 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2828 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2829 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2830 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2831 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2832 ] = { 5'd10,	5'd15,	5'd2,	5'd9};
	rom[ 2833 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2834 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2835 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2836 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2837 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2838 ] = { 5'd8,	5'd14,	5'd4,	5'd5};
	rom[ 2839 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2840 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2841 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2842 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2843 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2844 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2845 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2846 ] = { 5'd0,	5'd7,	5'd12,	5'd3};
	rom[ 2847 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2848 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2849 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2850 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2851 ] = { 5'd12,	5'd22,	5'd11,	5'd2};
	rom[ 2852 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2853 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2854 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2855 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2856 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2857 ] = { 5'd11,	5'd9,	5'd9,	5'd3};
	rom[ 2858 ] = { 5'd10,	5'd15,	5'd2,	5'd9};
	rom[ 2859 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2860 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2861 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2862 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2863 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2864 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2865 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2866 ] = { 5'd6,	5'd12,	5'd8,	5'd3};
	rom[ 2867 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2868 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2869 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2870 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2871 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2872 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2873 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2874 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2875 ] = { 5'd5,	5'd7,	5'd3,	5'd7};
	rom[ 2876 ] = { 5'd15,	5'd8,	5'd3,	5'd7};
	rom[ 2877 ] = { 5'd6,	5'd8,	5'd3,	5'd7};
	rom[ 2878 ] = { 5'd3,	5'd22,	5'd9,	5'd2};
	rom[ 2879 ] = { 5'd7,	5'd10,	5'd2,	5'd10};
	rom[ 2880 ] = { 5'd16,	5'd14,	5'd4,	5'd6};
	rom[ 2881 ] = { 5'd4,	5'd14,	5'd4,	5'd6};
	rom[ 2882 ] = { 5'd13,	5'd17,	5'd5,	5'd4};
	rom[ 2883 ] = { 5'd6,	5'd17,	5'd5,	5'd4};
	rom[ 2884 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2885 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2886 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2887 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2888 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2889 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2890 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2891 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2892 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2893 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2894 ] = { 5'd11,	5'd18,	5'd5,	5'd4};
	rom[ 2895 ] = { 5'd11,	5'd21,	5'd11,	5'd3};
	rom[ 2896 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2897 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2898 ] = { 5'd18,	5'd18,	5'd3,	5'd6};
	rom[ 2899 ] = { 5'd3,	5'd18,	5'd3,	5'd6};
	rom[ 2900 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2901 ] = { 5'd12,	5'd11,	5'd11,	5'd5};
	rom[ 2902 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2903 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2904 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2905 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2906 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2907 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2908 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2909 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2910 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2911 ] = { 5'd0,	5'd0,	5'd0,	5'd0};
	rom[ 2912 ] = { 5'd9,	5'd12,	5'd3,	5'd11};
	
	end
endmodule

module rect0_wieght_rom(
	input 				clk,
	input		[11:0]	addr,
	output reg	[14:0]	q    // x y w h 5bit*4
	);
	reg					[14:0]	rom [4095:0];
	//always @(posedge clk) q <= rom[addr];
	always @(posedge clk) q <= -4096;

endmodule

module rect1_wieght_rom(
	input 				clk,
	input		[11:0]	addr,
	output reg	[14:0]	q    // x y w h 5bit*4
	);
	reg					[14:0]	rom [4095:0];
	always @(posedge clk) q <= rom[addr];
	initial begin
	rom[ 0    ] = 12288; 
	rom[ 1    ] = 12288; 
	rom[ 2    ] = 12288; 
	rom[ 3    ] = 12288; 
	rom[ 4    ] = 8192; 
	rom[ 5    ] = 8192; 
	rom[ 6    ] = 8192; 
	rom[ 7    ] = 8192; 
	rom[ 8    ] = 8192; 
	rom[ 9    ] = 12288; 
	rom[ 10   ] = 12288; 
	rom[ 11   ] = 12288; 
	rom[ 12   ] = 12288; 
	rom[ 13   ] = 12288; 
	rom[ 14   ] = 8192; 
	rom[ 15   ] = 12288; 
	rom[ 16   ] = 12288; 
	rom[ 17   ] = 12288; 
	rom[ 18   ] = 12288; 
	rom[ 19   ] = 8192; 
	rom[ 20   ] = 12288; 
	rom[ 21   ] = 12288; 
	rom[ 22   ] = 12288; 
	rom[ 23   ] = 12288; 
	rom[ 24   ] = 8192; 
	rom[ 25   ] = 12288; 
	rom[ 26   ] = 8192; 
	rom[ 27   ] = 8192; 
	rom[ 28   ] = 12288; 
	rom[ 29   ] = 8192; 
	rom[ 30   ] = 12288; 
	rom[ 31   ] = 12288; 
	rom[ 32   ] = 8192; 
	rom[ 33   ] = 8192; 
	rom[ 34   ] = 12288; 
	rom[ 35   ] = 8192; 
	rom[ 36   ] = 12288; 
	rom[ 37   ] = 8192; 
	rom[ 38   ] = 8192; 
	rom[ 39   ] = 12288; 
	rom[ 40   ] = 8192; 
	rom[ 41   ] = 8192; 
	rom[ 42   ] = 12288; 
	rom[ 43   ] = 12288; 
	rom[ 44   ] = 8192; 
	rom[ 45   ] = 12288; 
	rom[ 46   ] = 8192; 
	rom[ 47   ] = 8192; 
	rom[ 48   ] = 8192; 
	rom[ 49   ] = 8192; 
	rom[ 50   ] = 8192; 
	rom[ 51   ] = 12288; 
	rom[ 52   ] = 12288; 
	rom[ 53   ] = 12288; 
	rom[ 54   ] = 12288; 
	rom[ 55   ] = 12288; 
	rom[ 56   ] = 8192; 
	rom[ 57   ] = 8192; 
	rom[ 58   ] = 8192; 
	rom[ 59   ] = 12288; 
	rom[ 60   ] = 12288; 
	rom[ 61   ] = 8192; 
	rom[ 62   ] = 8192; 
	rom[ 63   ] = 12288; 
	rom[ 64   ] = 8192; 
	rom[ 65   ] = 12288; 
	rom[ 66   ] = 12288; 
	rom[ 67   ] = 8192; 
	rom[ 68   ] = 8192; 
	rom[ 69   ] = 8192; 
	rom[ 70   ] = 8192; 
	rom[ 71   ] = 12288; 
	rom[ 72   ] = 12288; 
	rom[ 73   ] = 12288; 
	rom[ 74   ] = 12288; 
	rom[ 75   ] = 8192; 
	rom[ 76   ] = 8192; 
	rom[ 77   ] = 12288; 
	rom[ 78   ] = 12288; 
	rom[ 79   ] = 12288; 
	rom[ 80   ] = 12288; 
	rom[ 81   ] = 12288; 
	rom[ 82   ] = 12288; 
	rom[ 83   ] = 12288; 
	rom[ 84   ] = 12288; 
	rom[ 85   ] = 12288; 
	rom[ 86   ] = 12288; 
	rom[ 87   ] = 8192; 
	rom[ 88   ] = 12288; 
	rom[ 89   ] = 8192; 
	rom[ 90   ] = 12288; 
	rom[ 91   ] = 8192; 
	rom[ 92   ] = 8192; 
	rom[ 93   ] = 8192; 
	rom[ 94   ] = 8192; 
	rom[ 95   ] = 8192; 
	rom[ 96   ] = 8192; 
	rom[ 97   ] = 12288; 
	rom[ 98   ] = 8192; 
	rom[ 99   ] = 8192; 
	rom[ 100  ] = 12288; 
	rom[ 101  ] = 12288; 
	rom[ 102  ] = 8192; 
	rom[ 103  ] = 8192; 
	rom[ 104  ] = 8192; 
	rom[ 105  ] = 8192; 
	rom[ 106  ] = 8192; 
	rom[ 107  ] = 12288; 
	rom[ 108  ] = 8192; 
	rom[ 109  ] = 8192; 
	rom[ 110  ] = 8192; 
	rom[ 111  ] = 12288; 
	rom[ 112  ] = 12288; 
	rom[ 113  ] = 12288; 
	rom[ 114  ] = 12288; 
	rom[ 115  ] = 12288; 
	rom[ 116  ] = 8192; 
	rom[ 117  ] = 8192; 
	rom[ 118  ] = 8192; 
	rom[ 119  ] = 8192; 
	rom[ 120  ] = 8192; 
	rom[ 121  ] = 8192; 
	rom[ 122  ] = 8192; 
	rom[ 123  ] = 12288; 
	rom[ 124  ] = 8192; 
	rom[ 125  ] = 8192; 
	rom[ 126  ] = 8192; 
	rom[ 127  ] = 12288; 
	rom[ 128  ] = 8192; 
	rom[ 129  ] = 8192; 
	rom[ 130  ] = 8192; 
	rom[ 131  ] = 8192; 
	rom[ 132  ] = 12288; 
	rom[ 133  ] = 12288; 
	rom[ 134  ] = 12288; 
	rom[ 135  ] = 12288; 
	rom[ 136  ] = 12288; 
	rom[ 137  ] = 8192; 
	rom[ 138  ] = 12288; 
	rom[ 139  ] = 8192; 
	rom[ 140  ] = 12288; 
	rom[ 141  ] = 12288; 
	rom[ 142  ] = 12288; 
	rom[ 143  ] = 8192; 
	rom[ 144  ] = 8192; 
	rom[ 145  ] = 8192; 
	rom[ 146  ] = 8192; 
	rom[ 147  ] = 8192; 
	rom[ 148  ] = 12288; 
	rom[ 149  ] = 12288; 
	rom[ 150  ] = 12288; 
	rom[ 151  ] = 8192; 
	rom[ 152  ] = 8192; 
	rom[ 153  ] = 12288; 
	rom[ 154  ] = 12288; 
	rom[ 155  ] = 8192; 
	rom[ 156  ] = 8192; 
	rom[ 157  ] = 12288; 
	rom[ 158  ] = 8192; 
	rom[ 159  ] = 8192; 
	rom[ 160  ] = 8192; 
	rom[ 161  ] = 12288; 
	rom[ 162  ] = 8192; 
	rom[ 163  ] = 12288; 
	rom[ 164  ] = 8192; 
	rom[ 165  ] = 12288; 
	rom[ 166  ] = 12288; 
	rom[ 167  ] = 12288; 
	rom[ 168  ] = 12288; 
	rom[ 169  ] = 12288; 
	rom[ 170  ] = 12288; 
	rom[ 171  ] = 12288; 
	rom[ 172  ] = 8192; 
	rom[ 173  ] = 8192; 
	rom[ 174  ] = 8192; 
	rom[ 175  ] = 12288; 
	rom[ 176  ] = 8192; 
	rom[ 177  ] = 8192; 
	rom[ 178  ] = 8192; 
	rom[ 179  ] = 8192; 
	rom[ 180  ] = 8192; 
	rom[ 181  ] = 8192; 
	rom[ 182  ] = 8192; 
	rom[ 183  ] = 12288; 
	rom[ 184  ] = 12288; 
	rom[ 185  ] = 8192; 
	rom[ 186  ] = 12288; 
	rom[ 187  ] = 8192; 
	rom[ 188  ] = 12288; 
	rom[ 189  ] = 8192; 
	rom[ 190  ] = 8192; 
	rom[ 191  ] = 8192; 
	rom[ 192  ] = 8192; 
	rom[ 193  ] = 12288; 
	rom[ 194  ] = 12288; 
	rom[ 195  ] = 8192; 
	rom[ 196  ] = 8192; 
	rom[ 197  ] = 12288; 
	rom[ 198  ] = 8192; 
	rom[ 199  ] = 8192; 
	rom[ 200  ] = 12288; 
	rom[ 201  ] = 12288; 
	rom[ 202  ] = 8192; 
	rom[ 203  ] = 8192; 
	rom[ 204  ] = 12288; 
	rom[ 205  ] = 12288; 
	rom[ 206  ] = 8192; 
	rom[ 207  ] = 8192; 
	rom[ 208  ] = 12288; 
	rom[ 209  ] = 12288; 
	rom[ 210  ] = 8192; 
	rom[ 211  ] = 8192; 
	rom[ 212  ] = 12288; 
	rom[ 213  ] = 12288; 
	rom[ 214  ] = 12288; 
	rom[ 215  ] = 8192; 
	rom[ 216  ] = 12288; 
	rom[ 217  ] = 8192; 
	rom[ 218  ] = 8192; 
	rom[ 219  ] = 8192; 
	rom[ 220  ] = 12288; 
	rom[ 221  ] = 12288; 
	rom[ 222  ] = 12288; 
	rom[ 223  ] = 8192; 
	rom[ 224  ] = 8192; 
	rom[ 225  ] = 12288; 
	rom[ 226  ] = 12288; 
	rom[ 227  ] = 8192; 
	rom[ 228  ] = 12288; 
	rom[ 229  ] = 12288; 
	rom[ 230  ] = 8192; 
	rom[ 231  ] = 12288; 
	rom[ 232  ] = 12288; 
	rom[ 233  ] = 12288; 
	rom[ 234  ] = 8192; 
	rom[ 235  ] = 8192; 
	rom[ 236  ] = 8192; 
	rom[ 237  ] = 8192; 
	rom[ 238  ] = 12288; 
	rom[ 239  ] = 12288; 
	rom[ 240  ] = 8192; 
	rom[ 241  ] = 8192; 
	rom[ 242  ] = 8192; 
	rom[ 243  ] = 12288; 
	rom[ 244  ] = 12288; 
	rom[ 245  ] = 8192; 
	rom[ 246  ] = 8192; 
	rom[ 247  ] = 8192; 
	rom[ 248  ] = 8192; 
	rom[ 249  ] = 8192; 
	rom[ 250  ] = 12288; 
	rom[ 251  ] = 12288; 
	rom[ 252  ] = 12288; 
	rom[ 253  ] = 12288; 
	rom[ 254  ] = 8192; 
	rom[ 255  ] = 8192; 
	rom[ 256  ] = 12288; 
	rom[ 257  ] = 8192; 
	rom[ 258  ] = 12288; 
	rom[ 259  ] = 12288; 
	rom[ 260  ] = 12288; 
	rom[ 261  ] = 8192; 
	rom[ 262  ] = 8192; 
	rom[ 263  ] = 8192; 
	rom[ 264  ] = 8192; 
	rom[ 265  ] = 12288; 
	rom[ 266  ] = 8192; 
	rom[ 267  ] = 12288; 
	rom[ 268  ] = 8192; 
	rom[ 269  ] = 8192; 
	rom[ 270  ] = 12288; 
	rom[ 271  ] = 12288; 
	rom[ 272  ] = 8192; 
	rom[ 273  ] = 12288; 
	rom[ 274  ] = 12288; 
	rom[ 275  ] = 12288; 
	rom[ 276  ] = 8192; 
	rom[ 277  ] = 12288; 
	rom[ 278  ] = 8192; 
	rom[ 279  ] = 8192; 
	rom[ 280  ] = 8192; 
	rom[ 281  ] = 8192; 
	rom[ 282  ] = 12288; 
	rom[ 283  ] = 12288; 
	rom[ 284  ] = 12288; 
	rom[ 285  ] = 12288; 
	rom[ 286  ] = 8192; 
	rom[ 287  ] = 8192; 
	rom[ 288  ] = 8192; 
	rom[ 289  ] = 12288; 
	rom[ 290  ] = 12288; 
	rom[ 291  ] = 8192; 
	rom[ 292  ] = 8192; 
	rom[ 293  ] = 8192; 
	rom[ 294  ] = 12288; 
	rom[ 295  ] = 8192; 
	rom[ 296  ] = 12288; 
	rom[ 297  ] = 12288; 
	rom[ 298  ] = 8192; 
	rom[ 299  ] = 12288; 
	rom[ 300  ] = 12288; 
	rom[ 301  ] = 12288; 
	rom[ 302  ] = 12288; 
	rom[ 303  ] = 12288; 
	rom[ 304  ] = 8192; 
	rom[ 305  ] = 8192; 
	rom[ 306  ] = 8192; 
	rom[ 307  ] = 8192; 
	rom[ 308  ] = 8192; 
	rom[ 309  ] = 12288; 
	rom[ 310  ] = 12288; 
	rom[ 311  ] = 12288; 
	rom[ 312  ] = 12288; 
	rom[ 313  ] = 12288; 
	rom[ 314  ] = 12288; 
	rom[ 315  ] = 12288; 
	rom[ 316  ] = 8192; 
	rom[ 317  ] = 8192; 
	rom[ 318  ] = 8192; 
	rom[ 319  ] = 8192; 
	rom[ 320  ] = 8192; 
	rom[ 321  ] = 12288; 
	rom[ 322  ] = 12288; 
	rom[ 323  ] = 12288; 
	rom[ 324  ] = 12288; 
	rom[ 325  ] = 12288; 
	rom[ 326  ] = 12288; 
	rom[ 327  ] = 8192; 
	rom[ 328  ] = 8192; 
	rom[ 329  ] = 8192; 
	rom[ 330  ] = 12288; 
	rom[ 331  ] = 8192; 
	rom[ 332  ] = 12288; 
	rom[ 333  ] = 12288; 
	rom[ 334  ] = 8192; 
	rom[ 335  ] = 12288; 
	rom[ 336  ] = 8192; 
	rom[ 337  ] = 8192; 
	rom[ 338  ] = 12288; 
	rom[ 339  ] = 12288; 
	rom[ 340  ] = 12288; 
	rom[ 341  ] = 12288; 
	rom[ 342  ] = 8192; 
	rom[ 343  ] = 12288; 
	rom[ 344  ] = 12288; 
	rom[ 345  ] = 12288; 
	rom[ 346  ] = 12288; 
	rom[ 347  ] = 12288; 
	rom[ 348  ] = 12288; 
	rom[ 349  ] = 8192; 
	rom[ 350  ] = 12288; 
	rom[ 351  ] = 8192; 
	rom[ 352  ] = 12288; 
	rom[ 353  ] = 8192; 
	rom[ 354  ] = 8192; 
	rom[ 355  ] = 8192; 
	rom[ 356  ] = 12288; 
	rom[ 357  ] = 12288; 
	rom[ 358  ] = 12288; 
	rom[ 359  ] = 8192; 
	rom[ 360  ] = 8192; 
	rom[ 361  ] = 8192; 
	rom[ 362  ] = 8192; 
	rom[ 363  ] = 8192; 
	rom[ 364  ] = 12288; 
	rom[ 365  ] = 12288; 
	rom[ 366  ] = 8192; 
	rom[ 367  ] = 8192; 
	rom[ 368  ] = 12288; 
	rom[ 369  ] = 12288; 
	rom[ 370  ] = 12288; 
	rom[ 371  ] = 12288; 
	rom[ 372  ] = 12288; 
	rom[ 373  ] = 8192; 
	rom[ 374  ] = 8192; 
	rom[ 375  ] = 8192; 
	rom[ 376  ] = 12288; 
	rom[ 377  ] = 8192; 
	rom[ 378  ] = 8192; 
	rom[ 379  ] = 8192; 
	rom[ 380  ] = 12288; 
	rom[ 381  ] = 12288; 
	rom[ 382  ] = 12288; 
	rom[ 383  ] = 12288; 
	rom[ 384  ] = 8192; 
	rom[ 385  ] = 12288; 
	rom[ 386  ] = 12288; 
	rom[ 387  ] = 12288; 
	rom[ 388  ] = 12288; 
	rom[ 389  ] = 12288; 
	rom[ 390  ] = 12288; 
	rom[ 391  ] = 12288; 
	rom[ 392  ] = 8192; 
	rom[ 393  ] = 12288; 
	rom[ 394  ] = 12288; 
	rom[ 395  ] = 12288; 
	rom[ 396  ] = 12288; 
	rom[ 397  ] = 12288; 
	rom[ 398  ] = 8192; 
	rom[ 399  ] = 12288; 
	rom[ 400  ] = 12288; 
	rom[ 401  ] = 12288; 
	rom[ 402  ] = 12288; 
	rom[ 403  ] = 8192; 
	rom[ 404  ] = 8192; 
	rom[ 405  ] = 12288; 
	rom[ 406  ] = 12288; 
	rom[ 407  ] = 12288; 
	rom[ 408  ] = 12288; 
	rom[ 409  ] = 12288; 
	rom[ 410  ] = 8192; 
	rom[ 411  ] = 12288; 
	rom[ 412  ] = 8192; 
	rom[ 413  ] = 8192; 
	rom[ 414  ] = 8192; 
	rom[ 415  ] = 8192; 
	rom[ 416  ] = 8192; 
	rom[ 417  ] = 12288; 
	rom[ 418  ] = 12288; 
	rom[ 419  ] = 12288; 
	rom[ 420  ] = 12288; 
	rom[ 421  ] = 8192; 
	rom[ 422  ] = 8192; 
	rom[ 423  ] = 12288; 
	rom[ 424  ] = 12288; 
	rom[ 425  ] = 12288; 
	rom[ 426  ] = 8192; 
	rom[ 427  ] = 12288; 
	rom[ 428  ] = 12288; 
	rom[ 429  ] = 12288; 
	rom[ 430  ] = 12288; 
	rom[ 431  ] = 8192; 
	rom[ 432  ] = 8192; 
	rom[ 433  ] = 12288; 
	rom[ 434  ] = 12288; 
	rom[ 435  ] = 8192; 
	rom[ 436  ] = 8192; 
	rom[ 437  ] = 12288; 
	rom[ 438  ] = 8192; 
	rom[ 439  ] = 12288; 
	rom[ 440  ] = 12288; 
	rom[ 441  ] = 12288; 
	rom[ 442  ] = 12288; 
	rom[ 443  ] = 8192; 
	rom[ 444  ] = 8192; 
	rom[ 445  ] = 8192; 
	rom[ 446  ] = 8192; 
	rom[ 447  ] = 12288; 
	rom[ 448  ] = 8192; 
	rom[ 449  ] = 12288; 
	rom[ 450  ] = 12288; 
	rom[ 451  ] = 8192; 
	rom[ 452  ] = 8192; 
	rom[ 453  ] = 8192; 
	rom[ 454  ] = 8192; 
	rom[ 455  ] = 8192; 
	rom[ 456  ] = 8192; 
	rom[ 457  ] = 8192; 
	rom[ 458  ] = 12288; 
	rom[ 459  ] = 8192; 
	rom[ 460  ] = 8192; 
	rom[ 461  ] = 8192; 
	rom[ 462  ] = 12288; 
	rom[ 463  ] = 8192; 
	rom[ 464  ] = 8192; 
	rom[ 465  ] = 12288; 
	rom[ 466  ] = 8192; 
	rom[ 467  ] = 12288; 
	rom[ 468  ] = 12288; 
	rom[ 469  ] = 12288; 
	rom[ 470  ] = 8192; 
	rom[ 471  ] = 12288; 
	rom[ 472  ] = 12288; 
	rom[ 473  ] = 8192; 
	rom[ 474  ] = 8192; 
	rom[ 475  ] = 12288; 
	rom[ 476  ] = 12288; 
	rom[ 477  ] = 12288; 
	rom[ 478  ] = 8192; 
	rom[ 479  ] = 12288; 
	rom[ 480  ] = 12288; 
	rom[ 481  ] = 8192; 
	rom[ 482  ] = 8192; 
	rom[ 483  ] = 12288; 
	rom[ 484  ] = 12288; 
	rom[ 485  ] = 12288; 
	rom[ 486  ] = 12288; 
	rom[ 487  ] = 8192; 
	rom[ 488  ] = 8192; 
	rom[ 489  ] = 8192; 
	rom[ 490  ] = 8192; 
	rom[ 491  ] = 12288; 
	rom[ 492  ] = 12288; 
	rom[ 493  ] = 12288; 
	rom[ 494  ] = 12288; 
	rom[ 495  ] = 8192; 
	rom[ 496  ] = 8192; 
	rom[ 497  ] = 12288; 
	rom[ 498  ] = 12288; 
	rom[ 499  ] = 12288; 
	rom[ 500  ] = 12288; 
	rom[ 501  ] = 12288; 
	rom[ 502  ] = 12288; 
	rom[ 503  ] = 12288; 
	rom[ 504  ] = 12288; 
	rom[ 505  ] = 8192; 
	rom[ 506  ] = 12288; 
	rom[ 507  ] = 12288; 
	rom[ 508  ] = 12288; 
	rom[ 509  ] = 8192; 
	rom[ 510  ] = 12288; 
	rom[ 511  ] = 12288; 
	rom[ 512  ] = 12288; 
	rom[ 513  ] = 12288; 
	rom[ 514  ] = 12288; 
	rom[ 515  ] = 12288; 
	rom[ 516  ] = 12288; 
	rom[ 517  ] = 8192; 
	rom[ 518  ] = 12288; 
	rom[ 519  ] = 12288; 
	rom[ 520  ] = 8192; 
	rom[ 521  ] = 8192; 
	rom[ 522  ] = 8192; 
	rom[ 523  ] = 8192; 
	rom[ 524  ] = 8192; 
	rom[ 525  ] = 8192; 
	rom[ 526  ] = 12288; 
	rom[ 527  ] = 12288; 
	rom[ 528  ] = 12288; 
	rom[ 529  ] = 8192; 
	rom[ 530  ] = 12288; 
	rom[ 531  ] = 8192; 
	rom[ 532  ] = 12288; 
	rom[ 533  ] = 12288; 
	rom[ 534  ] = 12288; 
	rom[ 535  ] = 12288; 
	rom[ 536  ] = 12288; 
	rom[ 537  ] = 8192; 
	rom[ 538  ] = 8192; 
	rom[ 539  ] = 8192; 
	rom[ 540  ] = 8192; 
	rom[ 541  ] = 12288; 
	rom[ 542  ] = 8192; 
	rom[ 543  ] = 8192; 
	rom[ 544  ] = 12288; 
	rom[ 545  ] = 12288; 
	rom[ 546  ] = 8192; 
	rom[ 547  ] = 12288; 
	rom[ 548  ] = 8192; 
	rom[ 549  ] = 8192; 
	rom[ 550  ] = 8192; 
	rom[ 551  ] = 12288; 
	rom[ 552  ] = 8192; 
	rom[ 553  ] = 8192; 
	rom[ 554  ] = 8192; 
	rom[ 555  ] = 12288; 
	rom[ 556  ] = 12288; 
	rom[ 557  ] = 12288; 
	rom[ 558  ] = 12288; 
	rom[ 559  ] = 8192; 
	rom[ 560  ] = 12288; 
	rom[ 561  ] = 12288; 
	rom[ 562  ] = 12288; 
	rom[ 563  ] = 12288; 
	rom[ 564  ] = 8192; 
	rom[ 565  ] = 8192; 
	rom[ 566  ] = 8192; 
	rom[ 567  ] = 8192; 
	rom[ 568  ] = 12288; 
	rom[ 569  ] = 12288; 
	rom[ 570  ] = 12288; 
	rom[ 571  ] = 12288; 
	rom[ 572  ] = 8192; 
	rom[ 573  ] = 12288; 
	rom[ 574  ] = 8192; 
	rom[ 575  ] = 8192; 
	rom[ 576  ] = 12288; 
	rom[ 577  ] = 12288; 
	rom[ 578  ] = 12288; 
	rom[ 579  ] = 12288; 
	rom[ 580  ] = 12288; 
	rom[ 581  ] = 12288; 
	rom[ 582  ] = 12288; 
	rom[ 583  ] = 12288; 
	rom[ 584  ] = 8192; 
	rom[ 585  ] = 12288; 
	rom[ 586  ] = 12288; 
	rom[ 587  ] = 8192; 
	rom[ 588  ] = 8192; 
	rom[ 589  ] = 12288; 
	rom[ 590  ] = 12288; 
	rom[ 591  ] = 8192; 
	rom[ 592  ] = 8192; 
	rom[ 593  ] = 12288; 
	rom[ 594  ] = 8192; 
	rom[ 595  ] = 8192; 
	rom[ 596  ] = 12288; 
	rom[ 597  ] = 12288; 
	rom[ 598  ] = 8192; 
	rom[ 599  ] = 12288; 
	rom[ 600  ] = 8192; 
	rom[ 601  ] = 8192; 
	rom[ 602  ] = 8192; 
	rom[ 603  ] = 8192; 
	rom[ 604  ] = 12288; 
	rom[ 605  ] = 12288; 
	rom[ 606  ] = 8192; 
	rom[ 607  ] = 8192; 
	rom[ 608  ] = 12288; 
	rom[ 609  ] = 8192; 
	rom[ 610  ] = 12288; 
	rom[ 611  ] = 8192; 
	rom[ 612  ] = 8192; 
	rom[ 613  ] = 12288; 
	rom[ 614  ] = 8192; 
	rom[ 615  ] = 12288; 
	rom[ 616  ] = 12288; 
	rom[ 617  ] = 12288; 
	rom[ 618  ] = 12288; 
	rom[ 619  ] = 12288; 
	rom[ 620  ] = 8192; 
	rom[ 621  ] = 12288; 
	rom[ 622  ] = 8192; 
	rom[ 623  ] = 8192; 
	rom[ 624  ] = 8192; 
	rom[ 625  ] = 8192; 
	rom[ 626  ] = 8192; 
	rom[ 627  ] = 8192; 
	rom[ 628  ] = 12288; 
	rom[ 629  ] = 8192; 
	rom[ 630  ] = 8192; 
	rom[ 631  ] = 8192; 
	rom[ 632  ] = 12288; 
	rom[ 633  ] = 8192; 
	rom[ 634  ] = 12288; 
	rom[ 635  ] = 12288; 
	rom[ 636  ] = 12288; 
	rom[ 637  ] = 8192; 
	rom[ 638  ] = 12288; 
	rom[ 639  ] = 8192; 
	rom[ 640  ] = 12288; 
	rom[ 641  ] = 12288; 
	rom[ 642  ] = 12288; 
	rom[ 643  ] = 12288; 
	rom[ 644  ] = 8192; 
	rom[ 645  ] = 12288; 
	rom[ 646  ] = 12288; 
	rom[ 647  ] = 12288; 
	rom[ 648  ] = 8192; 
	rom[ 649  ] = 12288; 
	rom[ 650  ] = 12288; 
	rom[ 651  ] = 12288; 
	rom[ 652  ] = 12288; 
	rom[ 653  ] = 12288; 
	rom[ 654  ] = 12288; 
	rom[ 655  ] = 8192; 
	rom[ 656  ] = 12288; 
	rom[ 657  ] = 12288; 
	rom[ 658  ] = 12288; 
	rom[ 659  ] = 8192; 
	rom[ 660  ] = 12288; 
	rom[ 661  ] = 12288; 
	rom[ 662  ] = 12288; 
	rom[ 663  ] = 8192; 
	rom[ 664  ] = 8192; 
	rom[ 665  ] = 8192; 
	rom[ 666  ] = 8192; 
	rom[ 667  ] = 8192; 
	rom[ 668  ] = 12288; 
	rom[ 669  ] = 8192; 
	rom[ 670  ] = 8192; 
	rom[ 671  ] = 12288; 
	rom[ 672  ] = 12288; 
	rom[ 673  ] = 8192; 
	rom[ 674  ] = 8192; 
	rom[ 675  ] = 8192; 
	rom[ 676  ] = 12288; 
	rom[ 677  ] = 12288; 
	rom[ 678  ] = 8192; 
	rom[ 679  ] = 8192; 
	rom[ 680  ] = 8192; 
	rom[ 681  ] = 8192; 
	rom[ 682  ] = 8192; 
	rom[ 683  ] = 8192; 
	rom[ 684  ] = 8192; 
	rom[ 685  ] = 12288; 
	rom[ 686  ] = 8192; 
	rom[ 687  ] = 12288; 
	rom[ 688  ] = 12288; 
	rom[ 689  ] = 12288; 
	rom[ 690  ] = 8192; 
	rom[ 691  ] = 8192; 
	rom[ 692  ] = 12288; 
	rom[ 693  ] = 12288; 
	rom[ 694  ] = 8192; 
	rom[ 695  ] = 8192; 
	rom[ 696  ] = 8192; 
	rom[ 697  ] = 12288; 
	rom[ 698  ] = 12288; 
	rom[ 699  ] = 8192; 
	rom[ 700  ] = 8192; 
	rom[ 701  ] = 8192; 
	rom[ 702  ] = 12288; 
	rom[ 703  ] = 8192; 
	rom[ 704  ] = 8192; 
	rom[ 705  ] = 8192; 
	rom[ 706  ] = 8192; 
	rom[ 707  ] = 12288; 
	rom[ 708  ] = 12288; 
	rom[ 709  ] = 8192; 
	rom[ 710  ] = 8192; 
	rom[ 711  ] = 12288; 
	rom[ 712  ] = 12288; 
	rom[ 713  ] = 8192; 
	rom[ 714  ] = 8192; 
	rom[ 715  ] = 8192; 
	rom[ 716  ] = 12288; 
	rom[ 717  ] = 8192; 
	rom[ 718  ] = 8192; 
	rom[ 719  ] = 8192; 
	rom[ 720  ] = 12288; 
	rom[ 721  ] = 8192; 
	rom[ 722  ] = 8192; 
	rom[ 723  ] = 12288; 
	rom[ 724  ] = 8192; 
	rom[ 725  ] = 8192; 
	rom[ 726  ] = 8192; 
	rom[ 727  ] = 8192; 
	rom[ 728  ] = 8192; 
	rom[ 729  ] = 12288; 
	rom[ 730  ] = 12288; 
	rom[ 731  ] = 12288; 
	rom[ 732  ] = 12288; 
	rom[ 733  ] = 12288; 
	rom[ 734  ] = 12288; 
	rom[ 735  ] = 12288; 
	rom[ 736  ] = 12288; 
	rom[ 737  ] = 12288; 
	rom[ 738  ] = 12288; 
	rom[ 739  ] = 8192; 
	rom[ 740  ] = 8192; 
	rom[ 741  ] = 8192; 
	rom[ 742  ] = 8192; 
	rom[ 743  ] = 8192; 
	rom[ 744  ] = 12288; 
	rom[ 745  ] = 8192; 
	rom[ 746  ] = 12288; 
	rom[ 747  ] = 12288; 
	rom[ 748  ] = 12288; 
	rom[ 749  ] = 8192; 
	rom[ 750  ] = 8192; 
	rom[ 751  ] = 8192; 
	rom[ 752  ] = 8192; 
	rom[ 753  ] = 8192; 
	rom[ 754  ] = 12288; 
	rom[ 755  ] = 12288; 
	rom[ 756  ] = 8192; 
	rom[ 757  ] = 8192; 
	rom[ 758  ] = 8192; 
	rom[ 759  ] = 12288; 
	rom[ 760  ] = 12288; 
	rom[ 761  ] = 8192; 
	rom[ 762  ] = 12288; 
	rom[ 763  ] = 12288; 
	rom[ 764  ] = 8192; 
	rom[ 765  ] = 8192; 
	rom[ 766  ] = 8192; 
	rom[ 767  ] = 12288; 
	rom[ 768  ] = 12288; 
	rom[ 769  ] = 12288; 
	rom[ 770  ] = 8192; 
	rom[ 771  ] = 12288; 
	rom[ 772  ] = 12288; 
	rom[ 773  ] = 8192; 
	rom[ 774  ] = 12288; 
	rom[ 775  ] = 8192; 
	rom[ 776  ] = 8192; 
	rom[ 777  ] = 8192; 
	rom[ 778  ] = 8192; 
	rom[ 779  ] = 12288; 
	rom[ 780  ] = 8192; 
	rom[ 781  ] = 8192; 
	rom[ 782  ] = 8192; 
	rom[ 783  ] = 8192; 
	rom[ 784  ] = 8192; 
	rom[ 785  ] = 12288; 
	rom[ 786  ] = 8192; 
	rom[ 787  ] = 12288; 
	rom[ 788  ] = 12288; 
	rom[ 789  ] = 12288; 
	rom[ 790  ] = 12288; 
	rom[ 791  ] = 12288; 
	rom[ 792  ] = 12288; 
	rom[ 793  ] = 8192; 
	rom[ 794  ] = 8192; 
	rom[ 795  ] = 12288; 
	rom[ 796  ] = 12288; 
	rom[ 797  ] = 12288; 
	rom[ 798  ] = 8192; 
	rom[ 799  ] = 12288; 
	rom[ 800  ] = 8192; 
	rom[ 801  ] = 8192; 
	rom[ 802  ] = 12288; 
	rom[ 803  ] = 8192; 
	rom[ 804  ] = 8192; 
	rom[ 805  ] = 12288; 
	rom[ 806  ] = 12288; 
	rom[ 807  ] = 8192; 
	rom[ 808  ] = 12288; 
	rom[ 809  ] = 8192; 
	rom[ 810  ] = 8192; 
	rom[ 811  ] = 12288; 
	rom[ 812  ] = 8192; 
	rom[ 813  ] = 12288; 
	rom[ 814  ] = 12288; 
	rom[ 815  ] = 8192; 
	rom[ 816  ] = 8192; 
	rom[ 817  ] = 8192; 
	rom[ 818  ] = 12288; 
	rom[ 819  ] = 8192; 
	rom[ 820  ] = 12288; 
	rom[ 821  ] = 12288; 
	rom[ 822  ] = 12288; 
	rom[ 823  ] = 12288; 
	rom[ 824  ] = 8192; 
	rom[ 825  ] = 8192; 
	rom[ 826  ] = 12288; 
	rom[ 827  ] = 12288; 
	rom[ 828  ] = 8192; 
	rom[ 829  ] = 12288; 
	rom[ 830  ] = 12288; 
	rom[ 831  ] = 8192; 
	rom[ 832  ] = 12288; 
	rom[ 833  ] = 8192; 
	rom[ 834  ] = 12288; 
	rom[ 835  ] = 12288; 
	rom[ 836  ] = 12288; 
	rom[ 837  ] = 12288; 
	rom[ 838  ] = 12288; 
	rom[ 839  ] = 12288; 
	rom[ 840  ] = 12288; 
	rom[ 841  ] = 12288; 
	rom[ 842  ] = 8192; 
	rom[ 843  ] = 8192; 
	rom[ 844  ] = 8192; 
	rom[ 845  ] = 12288; 
	rom[ 846  ] = 12288; 
	rom[ 847  ] = 12288; 
	rom[ 848  ] = 12288; 
	rom[ 849  ] = 8192; 
	rom[ 850  ] = 8192; 
	rom[ 851  ] = 8192; 
	rom[ 852  ] = 12288; 
	rom[ 853  ] = 12288; 
	rom[ 854  ] = 12288; 
	rom[ 855  ] = 8192; 
	rom[ 856  ] = 8192; 
	rom[ 857  ] = 12288; 
	rom[ 858  ] = 12288; 
	rom[ 859  ] = 8192; 
	rom[ 860  ] = 12288; 
	rom[ 861  ] = 8192; 
	rom[ 862  ] = 8192; 
	rom[ 863  ] = 8192; 
	rom[ 864  ] = 8192; 
	rom[ 865  ] = 8192; 
	rom[ 866  ] = 8192; 
	rom[ 867  ] = 12288; 
	rom[ 868  ] = 8192; 
	rom[ 869  ] = 12288; 
	rom[ 870  ] = 8192; 
	rom[ 871  ] = 12288; 
	rom[ 872  ] = 8192; 
	rom[ 873  ] = 8192; 
	rom[ 874  ] = 8192; 
	rom[ 875  ] = 12288; 
	rom[ 876  ] = 8192; 
	rom[ 877  ] = 8192; 
	rom[ 878  ] = 12288; 
	rom[ 879  ] = 12288; 
	rom[ 880  ] = 12288; 
	rom[ 881  ] = 12288; 
	rom[ 882  ] = 12288; 
	rom[ 883  ] = 8192; 
	rom[ 884  ] = 12288; 
	rom[ 885  ] = 12288; 
	rom[ 886  ] = 12288; 
	rom[ 887  ] = 12288; 
	rom[ 888  ] = 12288; 
	rom[ 889  ] = 12288; 
	rom[ 890  ] = 12288; 
	rom[ 891  ] = 12288; 
	rom[ 892  ] = 8192; 
	rom[ 893  ] = 8192; 
	rom[ 894  ] = 8192; 
	rom[ 895  ] = 12288; 
	rom[ 896  ] = 8192; 
	rom[ 897  ] = 8192; 
	rom[ 898  ] = 12288; 
	rom[ 899  ] = 8192; 
	rom[ 900  ] = 8192; 
	rom[ 901  ] = 12288; 
	rom[ 902  ] = 8192; 
	rom[ 903  ] = 12288; 
	rom[ 904  ] = 8192; 
	rom[ 905  ] = 8192; 
	rom[ 906  ] = 8192; 
	rom[ 907  ] = 8192; 
	rom[ 908  ] = 8192; 
	rom[ 909  ] = 12288; 
	rom[ 910  ] = 12288; 
	rom[ 911  ] = 8192; 
	rom[ 912  ] = 8192; 
	rom[ 913  ] = 8192; 
	rom[ 914  ] = 12288; 
	rom[ 915  ] = 8192; 
	rom[ 916  ] = 12288; 
	rom[ 917  ] = 12288; 
	rom[ 918  ] = 12288; 
	rom[ 919  ] = 12288; 
	rom[ 920  ] = 8192; 
	rom[ 921  ] = 12288; 
	rom[ 922  ] = 8192; 
	rom[ 923  ] = 8192; 
	rom[ 924  ] = 12288; 
	rom[ 925  ] = 12288; 
	rom[ 926  ] = 12288; 
	rom[ 927  ] = 12288; 
	rom[ 928  ] = 12288; 
	rom[ 929  ] = 12288; 
	rom[ 930  ] = 12288; 
	rom[ 931  ] = 12288; 
	rom[ 932  ] = 12288; 
	rom[ 933  ] = 8192; 
	rom[ 934  ] = 8192; 
	rom[ 935  ] = 12288; 
	rom[ 936  ] = 12288; 
	rom[ 937  ] = 12288; 
	rom[ 938  ] = 12288; 
	rom[ 939  ] = 8192; 
	rom[ 940  ] = 8192; 
	rom[ 941  ] = 12288; 
	rom[ 942  ] = 12288; 
	rom[ 943  ] = 12288; 
	rom[ 944  ] = 12288; 
	rom[ 945  ] = 8192; 
	rom[ 946  ] = 8192; 
	rom[ 947  ] = 8192; 
	rom[ 948  ] = 12288; 
	rom[ 949  ] = 8192; 
	rom[ 950  ] = 8192; 
	rom[ 951  ] = 8192; 
	rom[ 952  ] = 12288; 
	rom[ 953  ] = 8192; 
	rom[ 954  ] = 8192; 
	rom[ 955  ] = 8192; 
	rom[ 956  ] = 8192; 
	rom[ 957  ] = 8192; 
	rom[ 958  ] = 12288; 
	rom[ 959  ] = 8192; 
	rom[ 960  ] = 8192; 
	rom[ 961  ] = 8192; 
	rom[ 962  ] = 8192; 
	rom[ 963  ] = 8192; 
	rom[ 964  ] = 8192; 
	rom[ 965  ] = 8192; 
	rom[ 966  ] = 8192; 
	rom[ 967  ] = 12288; 
	rom[ 968  ] = 8192; 
	rom[ 969  ] = 8192; 
	rom[ 970  ] = 12288; 
	rom[ 971  ] = 8192; 
	rom[ 972  ] = 8192; 
	rom[ 973  ] = 8192; 
	rom[ 974  ] = 12288; 
	rom[ 975  ] = 12288; 
	rom[ 976  ] = 12288; 
	rom[ 977  ] = 8192; 
	rom[ 978  ] = 8192; 
	rom[ 979  ] = 12288; 
	rom[ 980  ] = 8192; 
	rom[ 981  ] = 8192; 
	rom[ 982  ] = 8192; 
	rom[ 983  ] = 8192; 
	rom[ 984  ] = 8192; 
	rom[ 985  ] = 12288; 
	rom[ 986  ] = 8192; 
	rom[ 987  ] = 12288; 
	rom[ 988  ] = 8192; 
	rom[ 989  ] = 12288; 
	rom[ 990  ] = 8192; 
	rom[ 991  ] = 8192; 
	rom[ 992  ] = 12288; 
	rom[ 993  ] = 12288; 
	rom[ 994  ] = 8192; 
	rom[ 995  ] = 8192; 
	rom[ 996  ] = 12288; 
	rom[ 997  ] = 12288; 
	rom[ 998  ] = 8192; 
	rom[ 999  ] = 8192; 
	rom[ 1000 ] = 12288; 
	rom[ 1001 ] = 12288; 
	rom[ 1002 ] = 12288; 
	rom[ 1003 ] = 12288; 
	rom[ 1004 ] = 8192; 
	rom[ 1005 ] = 8192; 
	rom[ 1006 ] = 8192; 
	rom[ 1007 ] = 12288; 
	rom[ 1008 ] = 12288; 
	rom[ 1009 ] = 8192; 
	rom[ 1010 ] = 12288; 
	rom[ 1011 ] = 12288; 
	rom[ 1012 ] = 8192; 
	rom[ 1013 ] = 8192; 
	rom[ 1014 ] = 8192; 
	rom[ 1015 ] = 12288; 
	rom[ 1016 ] = 8192; 
	rom[ 1017 ] = 8192; 
	rom[ 1018 ] = 8192; 
	rom[ 1019 ] = 12288; 
	rom[ 1020 ] = 12288; 
	rom[ 1021 ] = 8192; 
	rom[ 1022 ] = 12288; 
	rom[ 1023 ] = 12288; 
	rom[ 1024 ] = 12288; 
	rom[ 1025 ] = 8192; 
	rom[ 1026 ] = 8192; 
	rom[ 1027 ] = 8192; 
	rom[ 1028 ] = 8192; 
	rom[ 1029 ] = 8192; 
	rom[ 1030 ] = 12288; 
	rom[ 1031 ] = 12288; 
	rom[ 1032 ] = 12288; 
	rom[ 1033 ] = 12288; 
	rom[ 1034 ] = 12288; 
	rom[ 1035 ] = 8192; 
	rom[ 1036 ] = 8192; 
	rom[ 1037 ] = 12288; 
	rom[ 1038 ] = 8192; 
	rom[ 1039 ] = 8192; 
	rom[ 1040 ] = 12288; 
	rom[ 1041 ] = 12288; 
	rom[ 1042 ] = 12288; 
	rom[ 1043 ] = 12288; 
	rom[ 1044 ] = 8192; 
	rom[ 1045 ] = 12288; 
	rom[ 1046 ] = 8192; 
	rom[ 1047 ] = 8192; 
	rom[ 1048 ] = 8192; 
	rom[ 1049 ] = 12288; 
	rom[ 1050 ] = 12288; 
	rom[ 1051 ] = 8192; 
	rom[ 1052 ] = 8192; 
	rom[ 1053 ] = 8192; 
	rom[ 1054 ] = 12288; 
	rom[ 1055 ] = 12288; 
	rom[ 1056 ] = 12288; 
	rom[ 1057 ] = 8192; 
	rom[ 1058 ] = 8192; 
	rom[ 1059 ] = 8192; 
	rom[ 1060 ] = 8192; 
	rom[ 1061 ] = 12288; 
	rom[ 1062 ] = 8192; 
	rom[ 1063 ] = 12288; 
	rom[ 1064 ] = 8192; 
	rom[ 1065 ] = 12288; 
	rom[ 1066 ] = 8192; 
	rom[ 1067 ] = 12288; 
	rom[ 1068 ] = 12288; 
	rom[ 1069 ] = 8192; 
	rom[ 1070 ] = 12288; 
	rom[ 1071 ] = 12288; 
	rom[ 1072 ] = 12288; 
	rom[ 1073 ] = 12288; 
	rom[ 1074 ] = 8192; 
	rom[ 1075 ] = 12288; 
	rom[ 1076 ] = 12288; 
	rom[ 1077 ] = 12288; 
	rom[ 1078 ] = 8192; 
	rom[ 1079 ] = 8192; 
	rom[ 1080 ] = 8192; 
	rom[ 1081 ] = 8192; 
	rom[ 1082 ] = 12288; 
	rom[ 1083 ] = 8192; 
	rom[ 1084 ] = 8192; 
	rom[ 1085 ] = 8192; 
	rom[ 1086 ] = 12288; 
	rom[ 1087 ] = 8192; 
	rom[ 1088 ] = 8192; 
	rom[ 1089 ] = 8192; 
	rom[ 1090 ] = 12288; 
	rom[ 1091 ] = 8192; 
	rom[ 1092 ] = 12288; 
	rom[ 1093 ] = 12288; 
	rom[ 1094 ] = 8192; 
	rom[ 1095 ] = 8192; 
	rom[ 1096 ] = 8192; 
	rom[ 1097 ] = 12288; 
	rom[ 1098 ] = 8192; 
	rom[ 1099 ] = 8192; 
	rom[ 1100 ] = 8192; 
	rom[ 1101 ] = 8192; 
	rom[ 1102 ] = 8192; 
	rom[ 1103 ] = 8192; 
	rom[ 1104 ] = 8192; 
	rom[ 1105 ] = 12288; 
	rom[ 1106 ] = 8192; 
	rom[ 1107 ] = 12288; 
	rom[ 1108 ] = 12288; 
	rom[ 1109 ] = 8192; 
	rom[ 1110 ] = 12288; 
	rom[ 1111 ] = 12288; 
	rom[ 1112 ] = 12288; 
	rom[ 1113 ] = 12288; 
	rom[ 1114 ] = 8192; 
	rom[ 1115 ] = 12288; 
	rom[ 1116 ] = 8192; 
	rom[ 1117 ] = 8192; 
	rom[ 1118 ] = 12288; 
	rom[ 1119 ] = 12288; 
	rom[ 1120 ] = 8192; 
	rom[ 1121 ] = 8192; 
	rom[ 1122 ] = 8192; 
	rom[ 1123 ] = 8192; 
	rom[ 1124 ] = 12288; 
	rom[ 1125 ] = 12288; 
	rom[ 1126 ] = 8192; 
	rom[ 1127 ] = 8192; 
	rom[ 1128 ] = 12288; 
	rom[ 1129 ] = 12288; 
	rom[ 1130 ] = 12288; 
	rom[ 1131 ] = 8192; 
	rom[ 1132 ] = 8192; 
	rom[ 1133 ] = 8192; 
	rom[ 1134 ] = 12288; 
	rom[ 1135 ] = 8192; 
	rom[ 1136 ] = 8192; 
	rom[ 1137 ] = 8192; 
	rom[ 1138 ] = 8192; 
	rom[ 1139 ] = 8192; 
	rom[ 1140 ] = 12288; 
	rom[ 1141 ] = 8192; 
	rom[ 1142 ] = 12288; 
	rom[ 1143 ] = 12288; 
	rom[ 1144 ] = 8192; 
	rom[ 1145 ] = 12288; 
	rom[ 1146 ] = 12288; 
	rom[ 1147 ] = 12288; 
	rom[ 1148 ] = 12288; 
	rom[ 1149 ] = 12288; 
	rom[ 1150 ] = 12288; 
	rom[ 1151 ] = 12288; 
	rom[ 1152 ] = 12288; 
	rom[ 1153 ] = 12288; 
	rom[ 1154 ] = 12288; 
	rom[ 1155 ] = 8192; 
	rom[ 1156 ] = 12288; 
	rom[ 1157 ] = 12288; 
	rom[ 1158 ] = 12288; 
	rom[ 1159 ] = 12288; 
	rom[ 1160 ] = 12288; 
	rom[ 1161 ] = 8192; 
	rom[ 1162 ] = 12288; 
	rom[ 1163 ] = 12288; 
	rom[ 1164 ] = 12288; 
	rom[ 1165 ] = 12288; 
	rom[ 1166 ] = 12288; 
	rom[ 1167 ] = 12288; 
	rom[ 1168 ] = 12288; 
	rom[ 1169 ] = 12288; 
	rom[ 1170 ] = 8192; 
	rom[ 1171 ] = 8192; 
	rom[ 1172 ] = 12288; 
	rom[ 1173 ] = 12288; 
	rom[ 1174 ] = 12288; 
	rom[ 1175 ] = 12288; 
	rom[ 1176 ] = 12288; 
	rom[ 1177 ] = 8192; 
	rom[ 1178 ] = 8192; 
	rom[ 1179 ] = 8192; 
	rom[ 1180 ] = 8192; 
	rom[ 1181 ] = 8192; 
	rom[ 1182 ] = 12288; 
	rom[ 1183 ] = 12288; 
	rom[ 1184 ] = 8192; 
	rom[ 1185 ] = 12288; 
	rom[ 1186 ] = 12288; 
	rom[ 1187 ] = 8192; 
	rom[ 1188 ] = 8192; 
	rom[ 1189 ] = 12288; 
	rom[ 1190 ] = 8192; 
	rom[ 1191 ] = 8192; 
	rom[ 1192 ] = 8192; 
	rom[ 1193 ] = 12288; 
	rom[ 1194 ] = 12288; 
	rom[ 1195 ] = 12288; 
	rom[ 1196 ] = 12288; 
	rom[ 1197 ] = 12288; 
	rom[ 1198 ] = 12288; 
	rom[ 1199 ] = 8192; 
	rom[ 1200 ] = 8192; 
	rom[ 1201 ] = 8192; 
	rom[ 1202 ] = 12288; 
	rom[ 1203 ] = 8192; 
	rom[ 1204 ] = 12288; 
	rom[ 1205 ] = 12288; 
	rom[ 1206 ] = 12288; 
	rom[ 1207 ] = 12288; 
	rom[ 1208 ] = 12288; 
	rom[ 1209 ] = 8192; 
	rom[ 1210 ] = 8192; 
	rom[ 1211 ] = 8192; 
	rom[ 1212 ] = 8192; 
	rom[ 1213 ] = 12288; 
	rom[ 1214 ] = 12288; 
	rom[ 1215 ] = 12288; 
	rom[ 1216 ] = 12288; 
	rom[ 1217 ] = 12288; 
	rom[ 1218 ] = 12288; 
	rom[ 1219 ] = 12288; 
	rom[ 1220 ] = 12288; 
	rom[ 1221 ] = 8192; 
	rom[ 1222 ] = 12288; 
	rom[ 1223 ] = 12288; 
	rom[ 1224 ] = 12288; 
	rom[ 1225 ] = 12288; 
	rom[ 1226 ] = 8192; 
	rom[ 1227 ] = 8192; 
	rom[ 1228 ] = 12288; 
	rom[ 1229 ] = 8192; 
	rom[ 1230 ] = 12288; 
	rom[ 1231 ] = 8192; 
	rom[ 1232 ] = 12288; 
	rom[ 1233 ] = 8192; 
	rom[ 1234 ] = 8192; 
	rom[ 1235 ] = 8192; 
	rom[ 1236 ] = 12288; 
	rom[ 1237 ] = 8192; 
	rom[ 1238 ] = 8192; 
	rom[ 1239 ] = 12288; 
	rom[ 1240 ] = 8192; 
	rom[ 1241 ] = 8192; 
	rom[ 1242 ] = 8192; 
	rom[ 1243 ] = 8192; 
	rom[ 1244 ] = 8192; 
	rom[ 1245 ] = 12288; 
	rom[ 1246 ] = 12288; 
	rom[ 1247 ] = 12288; 
	rom[ 1248 ] = 8192; 
	rom[ 1249 ] = 12288; 
	rom[ 1250 ] = 8192; 
	rom[ 1251 ] = 8192; 
	rom[ 1252 ] = 12288; 
	rom[ 1253 ] = 8192; 
	rom[ 1254 ] = 12288; 
	rom[ 1255 ] = 12288; 
	rom[ 1256 ] = 8192; 
	rom[ 1257 ] = 12288; 
	rom[ 1258 ] = 12288; 
	rom[ 1259 ] = 12288; 
	rom[ 1260 ] = 12288; 
	rom[ 1261 ] = 8192; 
	rom[ 1262 ] = 8192; 
	rom[ 1263 ] = 8192; 
	rom[ 1264 ] = 8192; 
	rom[ 1265 ] = 8192; 
	rom[ 1266 ] = 8192; 
	rom[ 1267 ] = 12288; 
	rom[ 1268 ] = 12288; 
	rom[ 1269 ] = 12288; 
	rom[ 1270 ] = 12288; 
	rom[ 1271 ] = 8192; 
	rom[ 1272 ] = 8192; 
	rom[ 1273 ] = 12288; 
	rom[ 1274 ] = 12288; 
	rom[ 1275 ] = 12288; 
	rom[ 1276 ] = 12288; 
	rom[ 1277 ] = 12288; 
	rom[ 1278 ] = 12288; 
	rom[ 1279 ] = 12288; 
	rom[ 1280 ] = 12288; 
	rom[ 1281 ] = 12288; 
	rom[ 1282 ] = 12288; 
	rom[ 1283 ] = 12288; 
	rom[ 1284 ] = 12288; 
	rom[ 1285 ] = 12288; 
	rom[ 1286 ] = 12288; 
	rom[ 1287 ] = 12288; 
	rom[ 1288 ] = 12288; 
	rom[ 1289 ] = 8192; 
	rom[ 1290 ] = 12288; 
	rom[ 1291 ] = 8192; 
	rom[ 1292 ] = 8192; 
	rom[ 1293 ] = 8192; 
	rom[ 1294 ] = 12288; 
	rom[ 1295 ] = 8192; 
	rom[ 1296 ] = 8192; 
	rom[ 1297 ] = 8192; 
	rom[ 1298 ] = 8192; 
	rom[ 1299 ] = 8192; 
	rom[ 1300 ] = 8192; 
	rom[ 1301 ] = 8192; 
	rom[ 1302 ] = 8192; 
	rom[ 1303 ] = 8192; 
	rom[ 1304 ] = 8192; 
	rom[ 1305 ] = 8192; 
	rom[ 1306 ] = 8192; 
	rom[ 1307 ] = 8192; 
	rom[ 1308 ] = 8192; 
	rom[ 1309 ] = 12288; 
	rom[ 1310 ] = 12288; 
	rom[ 1311 ] = 12288; 
	rom[ 1312 ] = 8192; 
	rom[ 1313 ] = 12288; 
	rom[ 1314 ] = 12288; 
	rom[ 1315 ] = 8192; 
	rom[ 1316 ] = 12288; 
	rom[ 1317 ] = 12288; 
	rom[ 1318 ] = 12288; 
	rom[ 1319 ] = 8192; 
	rom[ 1320 ] = 12288; 
	rom[ 1321 ] = 12288; 
	rom[ 1322 ] = 12288; 
	rom[ 1323 ] = 12288; 
	rom[ 1324 ] = 8192; 
	rom[ 1325 ] = 8192; 
	rom[ 1326 ] = 8192; 
	rom[ 1327 ] = 8192; 
	rom[ 1328 ] = 12288; 
	rom[ 1329 ] = 8192; 
	rom[ 1330 ] = 8192; 
	rom[ 1331 ] = 12288; 
	rom[ 1332 ] = 12288; 
	rom[ 1333 ] = 12288; 
	rom[ 1334 ] = 12288; 
	rom[ 1335 ] = 8192; 
	rom[ 1336 ] = 8192; 
	rom[ 1337 ] = 8192; 
	rom[ 1338 ] = 8192; 
	rom[ 1339 ] = 8192; 
	rom[ 1340 ] = 8192; 
	rom[ 1341 ] = 12288; 
	rom[ 1342 ] = 12288; 
	rom[ 1343 ] = 8192; 
	rom[ 1344 ] = 8192; 
	rom[ 1345 ] = 12288; 
	rom[ 1346 ] = 8192; 
	rom[ 1347 ] = 12288; 
	rom[ 1348 ] = 8192; 
	rom[ 1349 ] = 12288; 
	rom[ 1350 ] = 12288; 
	rom[ 1351 ] = 12288; 
	rom[ 1352 ] = 12288; 
	rom[ 1353 ] = 8192; 
	rom[ 1354 ] = 8192; 
	rom[ 1355 ] = 8192; 
	rom[ 1356 ] = 12288; 
	rom[ 1357 ] = 8192; 
	rom[ 1358 ] = 8192; 
	rom[ 1359 ] = 12288; 
	rom[ 1360 ] = 8192; 
	rom[ 1361 ] = 12288; 
	rom[ 1362 ] = 12288; 
	rom[ 1363 ] = 12288; 
	rom[ 1364 ] = 8192; 
	rom[ 1365 ] = 12288; 
	rom[ 1366 ] = 12288; 
	rom[ 1367 ] = 12288; 
	rom[ 1368 ] = 12288; 
	rom[ 1369 ] = 8192; 
	rom[ 1370 ] = 8192; 
	rom[ 1371 ] = 8192; 
	rom[ 1372 ] = 8192; 
	rom[ 1373 ] = 8192; 
	rom[ 1374 ] = 12288; 
	rom[ 1375 ] = 12288; 
	rom[ 1376 ] = 12288; 
	rom[ 1377 ] = 8192; 
	rom[ 1378 ] = 12288; 
	rom[ 1379 ] = 12288; 
	rom[ 1380 ] = 8192; 
	rom[ 1381 ] = 8192; 
	rom[ 1382 ] = 8192; 
	rom[ 1383 ] = 8192; 
	rom[ 1384 ] = 8192; 
	rom[ 1385 ] = 12288; 
	rom[ 1386 ] = 12288; 
	rom[ 1387 ] = 12288; 
	rom[ 1388 ] = 12288; 
	rom[ 1389 ] = 8192; 
	rom[ 1390 ] = 8192; 
	rom[ 1391 ] = 8192; 
	rom[ 1392 ] = 8192; 
	rom[ 1393 ] = 8192; 
	rom[ 1394 ] = 8192; 
	rom[ 1395 ] = 12288; 
	rom[ 1396 ] = 12288; 
	rom[ 1397 ] = 12288; 
	rom[ 1398 ] = 8192; 
	rom[ 1399 ] = 8192; 
	rom[ 1400 ] = 8192; 
	rom[ 1401 ] = 12288; 
	rom[ 1402 ] = 8192; 
	rom[ 1403 ] = 12288; 
	rom[ 1404 ] = 8192; 
	rom[ 1405 ] = 12288; 
	rom[ 1406 ] = 8192; 
	rom[ 1407 ] = 8192; 
	rom[ 1408 ] = 8192; 
	rom[ 1409 ] = 8192; 
	rom[ 1410 ] = 12288; 
	rom[ 1411 ] = 8192; 
	rom[ 1412 ] = 8192; 
	rom[ 1413 ] = 8192; 
	rom[ 1414 ] = 12288; 
	rom[ 1415 ] = 8192; 
	rom[ 1416 ] = 8192; 
	rom[ 1417 ] = 8192; 
	rom[ 1418 ] = 8192; 
	rom[ 1419 ] = 8192; 
	rom[ 1420 ] = 12288; 
	rom[ 1421 ] = 8192; 
	rom[ 1422 ] = 8192; 
	rom[ 1423 ] = 8192; 
	rom[ 1424 ] = 8192; 
	rom[ 1425 ] = 8192; 
	rom[ 1426 ] = 12288; 
	rom[ 1427 ] = 8192; 
	rom[ 1428 ] = 12288; 
	rom[ 1429 ] = 12288; 
	rom[ 1430 ] = 12288; 
	rom[ 1431 ] = 12288; 
	rom[ 1432 ] = 12288; 
	rom[ 1433 ] = 12288; 
	rom[ 1434 ] = 12288; 
	rom[ 1435 ] = 12288; 
	rom[ 1436 ] = 8192; 
	rom[ 1437 ] = 8192; 
	rom[ 1438 ] = 8192; 
	rom[ 1439 ] = 8192; 
	rom[ 1440 ] = 12288; 
	rom[ 1441 ] = 12288; 
	rom[ 1442 ] = 12288; 
	rom[ 1443 ] = 12288; 
	rom[ 1444 ] = 12288; 
	rom[ 1445 ] = 12288; 
	rom[ 1446 ] = 12288; 
	rom[ 1447 ] = 12288; 
	rom[ 1448 ] = 8192; 
	rom[ 1449 ] = 12288; 
	rom[ 1450 ] = 12288; 
	rom[ 1451 ] = 8192; 
	rom[ 1452 ] = 8192; 
	rom[ 1453 ] = 12288; 
	rom[ 1454 ] = 8192; 
	rom[ 1455 ] = 12288; 
	rom[ 1456 ] = 12288; 
	rom[ 1457 ] = 12288; 
	rom[ 1458 ] = 12288; 
	rom[ 1459 ] = 8192; 
	rom[ 1460 ] = 8192; 
	rom[ 1461 ] = 8192; 
	rom[ 1462 ] = 8192; 
	rom[ 1463 ] = 12288; 
	rom[ 1464 ] = 8192; 
	rom[ 1465 ] = 12288; 
	rom[ 1466 ] = 12288; 
	rom[ 1467 ] = 8192; 
	rom[ 1468 ] = 8192; 
	rom[ 1469 ] = 8192; 
	rom[ 1470 ] = 8192; 
	rom[ 1471 ] = 8192; 
	rom[ 1472 ] = 8192; 
	rom[ 1473 ] = 8192; 
	rom[ 1474 ] = 8192; 
	rom[ 1475 ] = 8192; 
	rom[ 1476 ] = 12288; 
	rom[ 1477 ] = 12288; 
	rom[ 1478 ] = 12288; 
	rom[ 1479 ] = 8192; 
	rom[ 1480 ] = 12288; 
	rom[ 1481 ] = 8192; 
	rom[ 1482 ] = 8192; 
	rom[ 1483 ] = 8192; 
	rom[ 1484 ] = 8192; 
	rom[ 1485 ] = 8192; 
	rom[ 1486 ] = 12288; 
	rom[ 1487 ] = 8192; 
	rom[ 1488 ] = 8192; 
	rom[ 1489 ] = 8192; 
	rom[ 1490 ] = 8192; 
	rom[ 1491 ] = 8192; 
	rom[ 1492 ] = 8192; 
	rom[ 1493 ] = 8192; 
	rom[ 1494 ] = 12288; 
	rom[ 1495 ] = 12288; 
	rom[ 1496 ] = 8192; 
	rom[ 1497 ] = 8192; 
	rom[ 1498 ] = 12288; 
	rom[ 1499 ] = 12288; 
	rom[ 1500 ] = 8192; 
	rom[ 1501 ] = 12288; 
	rom[ 1502 ] = 8192; 
	rom[ 1503 ] = 8192; 
	rom[ 1504 ] = 8192; 
	rom[ 1505 ] = 8192; 
	rom[ 1506 ] = 8192; 
	rom[ 1507 ] = 12288; 
	rom[ 1508 ] = 8192; 
	rom[ 1509 ] = 8192; 
	rom[ 1510 ] = 8192; 
	rom[ 1511 ] = 8192; 
	rom[ 1512 ] = 12288; 
	rom[ 1513 ] = 8192; 
	rom[ 1514 ] = 12288; 
	rom[ 1515 ] = 8192; 
	rom[ 1516 ] = 12288; 
	rom[ 1517 ] = 8192; 
	rom[ 1518 ] = 12288; 
	rom[ 1519 ] = 12288; 
	rom[ 1520 ] = 8192; 
	rom[ 1521 ] = 8192; 
	rom[ 1522 ] = 12288; 
	rom[ 1523 ] = 12288; 
	rom[ 1524 ] = 8192; 
	rom[ 1525 ] = 12288; 
	rom[ 1526 ] = 12288; 
	rom[ 1527 ] = 8192; 
	rom[ 1528 ] = 12288; 
	rom[ 1529 ] = 12288; 
	rom[ 1530 ] = 8192; 
	rom[ 1531 ] = 12288; 
	rom[ 1532 ] = 8192; 
	rom[ 1533 ] = 12288; 
	rom[ 1534 ] = 12288; 
	rom[ 1535 ] = 8192; 
	rom[ 1536 ] = 8192; 
	rom[ 1537 ] = 12288; 
	rom[ 1538 ] = 8192; 
	rom[ 1539 ] = 12288; 
	rom[ 1540 ] = 12288; 
	rom[ 1541 ] = 8192; 
	rom[ 1542 ] = 8192; 
	rom[ 1543 ] = 12288; 
	rom[ 1544 ] = 8192; 
	rom[ 1545 ] = 8192; 
	rom[ 1546 ] = 8192; 
	rom[ 1547 ] = 8192; 
	rom[ 1548 ] = 8192; 
	rom[ 1549 ] = 8192; 
	rom[ 1550 ] = 8192; 
	rom[ 1551 ] = 8192; 
	rom[ 1552 ] = 12288; 
	rom[ 1553 ] = 8192; 
	rom[ 1554 ] = 8192; 
	rom[ 1555 ] = 8192; 
	rom[ 1556 ] = 8192; 
	rom[ 1557 ] = 12288; 
	rom[ 1558 ] = 8192; 
	rom[ 1559 ] = 8192; 
	rom[ 1560 ] = 12288; 
	rom[ 1561 ] = 12288; 
	rom[ 1562 ] = 12288; 
	rom[ 1563 ] = 12288; 
	rom[ 1564 ] = 8192; 
	rom[ 1565 ] = 8192; 
	rom[ 1566 ] = 8192; 
	rom[ 1567 ] = 8192; 
	rom[ 1568 ] = 12288; 
	rom[ 1569 ] = 8192; 
	rom[ 1570 ] = 8192; 
	rom[ 1571 ] = 8192; 
	rom[ 1572 ] = 8192; 
	rom[ 1573 ] = 12288; 
	rom[ 1574 ] = 12288; 
	rom[ 1575 ] = 12288; 
	rom[ 1576 ] = 8192; 
	rom[ 1577 ] = 8192; 
	rom[ 1578 ] = 12288; 
	rom[ 1579 ] = 12288; 
	rom[ 1580 ] = 12288; 
	rom[ 1581 ] = 8192; 
	rom[ 1582 ] = 8192; 
	rom[ 1583 ] = 8192; 
	rom[ 1584 ] = 8192; 
	rom[ 1585 ] = 12288; 
	rom[ 1586 ] = 12288; 
	rom[ 1587 ] = 12288; 
	rom[ 1588 ] = 12288; 
	rom[ 1589 ] = 12288; 
	rom[ 1590 ] = 12288; 
	rom[ 1591 ] = 12288; 
	rom[ 1592 ] = 12288; 
	rom[ 1593 ] = 12288; 
	rom[ 1594 ] = 12288; 
	rom[ 1595 ] = 12288; 
	rom[ 1596 ] = 8192; 
	rom[ 1597 ] = 8192; 
	rom[ 1598 ] = 12288; 
	rom[ 1599 ] = 12288; 
	rom[ 1600 ] = 8192; 
	rom[ 1601 ] = 8192; 
	rom[ 1602 ] = 12288; 
	rom[ 1603 ] = 12288; 
	rom[ 1604 ] = 12288; 
	rom[ 1605 ] = 8192; 
	rom[ 1606 ] = 12288; 
	rom[ 1607 ] = 8192; 
	rom[ 1608 ] = 12288; 
	rom[ 1609 ] = 8192; 
	rom[ 1610 ] = 8192; 
	rom[ 1611 ] = 8192; 
	rom[ 1612 ] = 8192; 
	rom[ 1613 ] = 12288; 
	rom[ 1614 ] = 8192; 
	rom[ 1615 ] = 8192; 
	rom[ 1616 ] = 8192; 
	rom[ 1617 ] = 12288; 
	rom[ 1618 ] = 12288; 
	rom[ 1619 ] = 12288; 
	rom[ 1620 ] = 12288; 
	rom[ 1621 ] = 8192; 
	rom[ 1622 ] = 8192; 
	rom[ 1623 ] = 8192; 
	rom[ 1624 ] = 12288; 
	rom[ 1625 ] = 8192; 
	rom[ 1626 ] = 12288; 
	rom[ 1627 ] = 8192; 
	rom[ 1628 ] = 12288; 
	rom[ 1629 ] = 8192; 
	rom[ 1630 ] = 8192; 
	rom[ 1631 ] = 12288; 
	rom[ 1632 ] = 12288; 
	rom[ 1633 ] = 12288; 
	rom[ 1634 ] = 8192; 
	rom[ 1635 ] = 8192; 
	rom[ 1636 ] = 8192; 
	rom[ 1637 ] = 12288; 
	rom[ 1638 ] = 12288; 
	rom[ 1639 ] = 8192; 
	rom[ 1640 ] = 8192; 
	rom[ 1641 ] = 8192; 
	rom[ 1642 ] = 8192; 
	rom[ 1643 ] = 12288; 
	rom[ 1644 ] = 8192; 
	rom[ 1645 ] = 8192; 
	rom[ 1646 ] = 8192; 
	rom[ 1647 ] = 8192; 
	rom[ 1648 ] = 8192; 
	rom[ 1649 ] = 8192; 
	rom[ 1650 ] = 8192; 
	rom[ 1651 ] = 8192; 
	rom[ 1652 ] = 8192; 
	rom[ 1653 ] = 8192; 
	rom[ 1654 ] = 12288; 
	rom[ 1655 ] = 12288; 
	rom[ 1656 ] = 12288; 
	rom[ 1657 ] = 8192; 
	rom[ 1658 ] = 8192; 
	rom[ 1659 ] = 8192; 
	rom[ 1660 ] = 8192; 
	rom[ 1661 ] = 8192; 
	rom[ 1662 ] = 8192; 
	rom[ 1663 ] = 12288; 
	rom[ 1664 ] = 12288; 
	rom[ 1665 ] = 12288; 
	rom[ 1666 ] = 8192; 
	rom[ 1667 ] = 12288; 
	rom[ 1668 ] = 8192; 
	rom[ 1669 ] = 8192; 
	rom[ 1670 ] = 8192; 
	rom[ 1671 ] = 8192; 
	rom[ 1672 ] = 12288; 
	rom[ 1673 ] = 12288; 
	rom[ 1674 ] = 8192; 
	rom[ 1675 ] = 8192; 
	rom[ 1676 ] = 8192; 
	rom[ 1677 ] = 8192; 
	rom[ 1678 ] = 12288; 
	rom[ 1679 ] = 12288; 
	rom[ 1680 ] = 8192; 
	rom[ 1681 ] = 8192; 
	rom[ 1682 ] = 8192; 
	rom[ 1683 ] = 8192; 
	rom[ 1684 ] = 8192; 
	rom[ 1685 ] = 8192; 
	rom[ 1686 ] = 8192; 
	rom[ 1687 ] = 12288; 
	rom[ 1688 ] = 12288; 
	rom[ 1689 ] = 12288; 
	rom[ 1690 ] = 12288; 
	rom[ 1691 ] = 12288; 
	rom[ 1692 ] = 8192; 
	rom[ 1693 ] = 8192; 
	rom[ 1694 ] = 12288; 
	rom[ 1695 ] = 12288; 
	rom[ 1696 ] = 12288; 
	rom[ 1697 ] = 12288; 
	rom[ 1698 ] = 12288; 
	rom[ 1699 ] = 8192; 
	rom[ 1700 ] = 12288; 
	rom[ 1701 ] = 12288; 
	rom[ 1702 ] = 8192; 
	rom[ 1703 ] = 8192; 
	rom[ 1704 ] = 8192; 
	rom[ 1705 ] = 12288; 
	rom[ 1706 ] = 12288; 
	rom[ 1707 ] = 8192; 
	rom[ 1708 ] = 12288; 
	rom[ 1709 ] = 8192; 
	rom[ 1710 ] = 12288; 
	rom[ 1711 ] = 12288; 
	rom[ 1712 ] = 12288; 
	rom[ 1713 ] = 8192; 
	rom[ 1714 ] = 8192; 
	rom[ 1715 ] = 12288; 
	rom[ 1716 ] = 12288; 
	rom[ 1717 ] = 8192; 
	rom[ 1718 ] = 8192; 
	rom[ 1719 ] = 12288; 
	rom[ 1720 ] = 8192; 
	rom[ 1721 ] = 8192; 
	rom[ 1722 ] = 8192; 
	rom[ 1723 ] = 12288; 
	rom[ 1724 ] = 12288; 
	rom[ 1725 ] = 8192; 
	rom[ 1726 ] = 8192; 
	rom[ 1727 ] = 8192; 
	rom[ 1728 ] = 12288; 
	rom[ 1729 ] = 12288; 
	rom[ 1730 ] = 12288; 
	rom[ 1731 ] = 8192; 
	rom[ 1732 ] = 8192; 
	rom[ 1733 ] = 8192; 
	rom[ 1734 ] = 12288; 
	rom[ 1735 ] = 8192; 
	rom[ 1736 ] = 12288; 
	rom[ 1737 ] = 12288; 
	rom[ 1738 ] = 12288; 
	rom[ 1739 ] = 12288; 
	rom[ 1740 ] = 12288; 
	rom[ 1741 ] = 12288; 
	rom[ 1742 ] = 12288; 
	rom[ 1743 ] = 12288; 
	rom[ 1744 ] = 12288; 
	rom[ 1745 ] = 12288; 
	rom[ 1746 ] = 12288; 
	rom[ 1747 ] = 12288; 
	rom[ 1748 ] = 8192; 
	rom[ 1749 ] = 12288; 
	rom[ 1750 ] = 8192; 
	rom[ 1751 ] = 8192; 
	rom[ 1752 ] = 12288; 
	rom[ 1753 ] = 8192; 
	rom[ 1754 ] = 12288; 
	rom[ 1755 ] = 8192; 
	rom[ 1756 ] = 12288; 
	rom[ 1757 ] = 8192; 
	rom[ 1758 ] = 8192; 
	rom[ 1759 ] = 12288; 
	rom[ 1760 ] = 8192; 
	rom[ 1761 ] = 12288; 
	rom[ 1762 ] = 8192; 
	rom[ 1763 ] = 8192; 
	rom[ 1764 ] = 8192; 
	rom[ 1765 ] = 12288; 
	rom[ 1766 ] = 8192; 
	rom[ 1767 ] = 8192; 
	rom[ 1768 ] = 8192; 
	rom[ 1769 ] = 8192; 
	rom[ 1770 ] = 12288; 
	rom[ 1771 ] = 12288; 
	rom[ 1772 ] = 12288; 
	rom[ 1773 ] = 12288; 
	rom[ 1774 ] = 8192; 
	rom[ 1775 ] = 8192; 
	rom[ 1776 ] = 8192; 
	rom[ 1777 ] = 8192; 
	rom[ 1778 ] = 8192; 
	rom[ 1779 ] = 12288; 
	rom[ 1780 ] = 12288; 
	rom[ 1781 ] = 8192; 
	rom[ 1782 ] = 12288; 
	rom[ 1783 ] = 12288; 
	rom[ 1784 ] = 8192; 
	rom[ 1785 ] = 12288; 
	rom[ 1786 ] = 8192; 
	rom[ 1787 ] = 12288; 
	rom[ 1788 ] = 8192; 
	rom[ 1789 ] = 8192; 
	rom[ 1790 ] = 8192; 
	rom[ 1791 ] = 8192; 
	rom[ 1792 ] = 12288; 
	rom[ 1793 ] = 8192; 
	rom[ 1794 ] = 8192; 
	rom[ 1795 ] = 8192; 
	rom[ 1796 ] = 12288; 
	rom[ 1797 ] = 12288; 
	rom[ 1798 ] = 12288; 
	rom[ 1799 ] = 12288; 
	rom[ 1800 ] = 8192; 
	rom[ 1801 ] = 12288; 
	rom[ 1802 ] = 8192; 
	rom[ 1803 ] = 8192; 
	rom[ 1804 ] = 12288; 
	rom[ 1805 ] = 8192; 
	rom[ 1806 ] = 8192; 
	rom[ 1807 ] = 8192; 
	rom[ 1808 ] = 8192; 
	rom[ 1809 ] = 12288; 
	rom[ 1810 ] = 8192; 
	rom[ 1811 ] = 12288; 
	rom[ 1812 ] = 12288; 
	rom[ 1813 ] = 8192; 
	rom[ 1814 ] = 12288; 
	rom[ 1815 ] = 8192; 
	rom[ 1816 ] = 8192; 
	rom[ 1817 ] = 12288; 
	rom[ 1818 ] = 8192; 
	rom[ 1819 ] = 12288; 
	rom[ 1820 ] = 8192; 
	rom[ 1821 ] = 8192; 
	rom[ 1822 ] = 12288; 
	rom[ 1823 ] = 12288; 
	rom[ 1824 ] = 12288; 
	rom[ 1825 ] = 8192; 
	rom[ 1826 ] = 12288; 
	rom[ 1827 ] = 12288; 
	rom[ 1828 ] = 12288; 
	rom[ 1829 ] = 12288; 
	rom[ 1830 ] = 8192; 
	rom[ 1831 ] = 12288; 
	rom[ 1832 ] = 12288; 
	rom[ 1833 ] = 8192; 
	rom[ 1834 ] = 12288; 
	rom[ 1835 ] = 12288; 
	rom[ 1836 ] = 12288; 
	rom[ 1837 ] = 8192; 
	rom[ 1838 ] = 8192; 
	rom[ 1839 ] = 12288; 
	rom[ 1840 ] = 8192; 
	rom[ 1841 ] = 8192; 
	rom[ 1842 ] = 8192; 
	rom[ 1843 ] = 8192; 
	rom[ 1844 ] = 12288; 
	rom[ 1845 ] = 8192; 
	rom[ 1846 ] = 12288; 
	rom[ 1847 ] = 12288; 
	rom[ 1848 ] = 12288; 
	rom[ 1849 ] = 12288; 
	rom[ 1850 ] = 12288; 
	rom[ 1851 ] = 12288; 
	rom[ 1852 ] = 12288; 
	rom[ 1853 ] = 12288; 
	rom[ 1854 ] = 12288; 
	rom[ 1855 ] = 12288; 
	rom[ 1856 ] = 8192; 
	rom[ 1857 ] = 12288; 
	rom[ 1858 ] = 12288; 
	rom[ 1859 ] = 12288; 
	rom[ 1860 ] = 12288; 
	rom[ 1861 ] = 12288; 
	rom[ 1862 ] = 8192; 
	rom[ 1863 ] = 12288; 
	rom[ 1864 ] = 12288; 
	rom[ 1865 ] = 12288; 
	rom[ 1866 ] = 8192; 
	rom[ 1867 ] = 12288; 
	rom[ 1868 ] = 12288; 
	rom[ 1869 ] = 12288; 
	rom[ 1870 ] = 12288; 
	rom[ 1871 ] = 12288; 
	rom[ 1872 ] = 8192; 
	rom[ 1873 ] = 8192; 
	rom[ 1874 ] = 8192; 
	rom[ 1875 ] = 8192; 
	rom[ 1876 ] = 8192; 
	rom[ 1877 ] = 8192; 
	rom[ 1878 ] = 8192; 
	rom[ 1879 ] = 12288; 
	rom[ 1880 ] = 8192; 
	rom[ 1881 ] = 12288; 
	rom[ 1882 ] = 12288; 
	rom[ 1883 ] = 8192; 
	rom[ 1884 ] = 8192; 
	rom[ 1885 ] = 8192; 
	rom[ 1886 ] = 8192; 
	rom[ 1887 ] = 12288; 
	rom[ 1888 ] = 12288; 
	rom[ 1889 ] = 12288; 
	rom[ 1890 ] = 12288; 
	rom[ 1891 ] = 12288; 
	rom[ 1892 ] = 8192; 
	rom[ 1893 ] = 8192; 
	rom[ 1894 ] = 8192; 
	rom[ 1895 ] = 12288; 
	rom[ 1896 ] = 12288; 
	rom[ 1897 ] = 12288; 
	rom[ 1898 ] = 12288; 
	rom[ 1899 ] = 8192; 
	rom[ 1900 ] = 8192; 
	rom[ 1901 ] = 8192; 
	rom[ 1902 ] = 12288; 
	rom[ 1903 ] = 12288; 
	rom[ 1904 ] = 12288; 
	rom[ 1905 ] = 12288; 
	rom[ 1906 ] = 12288; 
	rom[ 1907 ] = 12288; 
	rom[ 1908 ] = 12288; 
	rom[ 1909 ] = 12288; 
	rom[ 1910 ] = 12288; 
	rom[ 1911 ] = 8192; 
	rom[ 1912 ] = 12288; 
	rom[ 1913 ] = 8192; 
	rom[ 1914 ] = 8192; 
	rom[ 1915 ] = 8192; 
	rom[ 1916 ] = 8192; 
	rom[ 1917 ] = 8192; 
	rom[ 1918 ] = 12288; 
	rom[ 1919 ] = 12288; 
	rom[ 1920 ] = 8192; 
	rom[ 1921 ] = 8192; 
	rom[ 1922 ] = 8192; 
	rom[ 1923 ] = 8192; 
	rom[ 1924 ] = 8192; 
	rom[ 1925 ] = 12288; 
	rom[ 1926 ] = 12288; 
	rom[ 1927 ] = 12288; 
	rom[ 1928 ] = 12288; 
	rom[ 1929 ] = 8192; 
	rom[ 1930 ] = 12288; 
	rom[ 1931 ] = 12288; 
	rom[ 1932 ] = 8192; 
	rom[ 1933 ] = 12288; 
	rom[ 1934 ] = 8192; 
	rom[ 1935 ] = 12288; 
	rom[ 1936 ] = 12288; 
	rom[ 1937 ] = 12288; 
	rom[ 1938 ] = 12288; 
	rom[ 1939 ] = 12288; 
	rom[ 1940 ] = 8192; 
	rom[ 1941 ] = 8192; 
	rom[ 1942 ] = 8192; 
	rom[ 1943 ] = 8192; 
	rom[ 1944 ] = 12288; 
	rom[ 1945 ] = 12288; 
	rom[ 1946 ] = 8192; 
	rom[ 1947 ] = 8192; 
	rom[ 1948 ] = 12288; 
	rom[ 1949 ] = 8192; 
	rom[ 1950 ] = 8192; 
	rom[ 1951 ] = 8192; 
	rom[ 1952 ] = 12288; 
	rom[ 1953 ] = 12288; 
	rom[ 1954 ] = 12288; 
	rom[ 1955 ] = 8192; 
	rom[ 1956 ] = 8192; 
	rom[ 1957 ] = 12288; 
	rom[ 1958 ] = 8192; 
	rom[ 1959 ] = 12288; 
	rom[ 1960 ] = 8192; 
	rom[ 1961 ] = 12288; 
	rom[ 1962 ] = 8192; 
	rom[ 1963 ] = 8192; 
	rom[ 1964 ] = 12288; 
	rom[ 1965 ] = 8192; 
	rom[ 1966 ] = 12288; 
	rom[ 1967 ] = 8192; 
	rom[ 1968 ] = 12288; 
	rom[ 1969 ] = 8192; 
	rom[ 1970 ] = 12288; 
	rom[ 1971 ] = 8192; 
	rom[ 1972 ] = 8192; 
	rom[ 1973 ] = 12288; 
	rom[ 1974 ] = 12288; 
	rom[ 1975 ] = 8192; 
	rom[ 1976 ] = 8192; 
	rom[ 1977 ] = 8192; 
	rom[ 1978 ] = 8192; 
	rom[ 1979 ] = 12288; 
	rom[ 1980 ] = 12288; 
	rom[ 1981 ] = 12288; 
	rom[ 1982 ] = 12288; 
	rom[ 1983 ] = 12288; 
	rom[ 1984 ] = 8192; 
	rom[ 1985 ] = 8192; 
	rom[ 1986 ] = 8192; 
	rom[ 1987 ] = 8192; 
	rom[ 1988 ] = 12288; 
	rom[ 1989 ] = 8192; 
	rom[ 1990 ] = 12288; 
	rom[ 1991 ] = 12288; 
	rom[ 1992 ] = 8192; 
	rom[ 1993 ] = 8192; 
	rom[ 1994 ] = 12288; 
	rom[ 1995 ] = 12288; 
	rom[ 1996 ] = 8192; 
	rom[ 1997 ] = 8192; 
	rom[ 1998 ] = 8192; 
	rom[ 1999 ] = 12288; 
	rom[ 2000 ] = 8192; 
	rom[ 2001 ] = 8192; 
	rom[ 2002 ] = 12288; 
	rom[ 2003 ] = 8192; 
	rom[ 2004 ] = 8192; 
	rom[ 2005 ] = 8192; 
	rom[ 2006 ] = 12288; 
	rom[ 2007 ] = 8192; 
	rom[ 2008 ] = 12288; 
	rom[ 2009 ] = 8192; 
	rom[ 2010 ] = 12288; 
	rom[ 2011 ] = 8192; 
	rom[ 2012 ] = 12288; 
	rom[ 2013 ] = 12288; 
	rom[ 2014 ] = 8192; 
	rom[ 2015 ] = 8192; 
	rom[ 2016 ] = 12288; 
	rom[ 2017 ] = 8192; 
	rom[ 2018 ] = 8192; 
	rom[ 2019 ] = 8192; 
	rom[ 2020 ] = 8192; 
	rom[ 2021 ] = 8192; 
	rom[ 2022 ] = 12288; 
	rom[ 2023 ] = 8192; 
	rom[ 2024 ] = 12288; 
	rom[ 2025 ] = 8192; 
	rom[ 2026 ] = 12288; 
	rom[ 2027 ] = 12288; 
	rom[ 2028 ] = 12288; 
	rom[ 2029 ] = 12288; 
	rom[ 2030 ] = 12288; 
	rom[ 2031 ] = 12288; 
	rom[ 2032 ] = 12288; 
	rom[ 2033 ] = 8192; 
	rom[ 2034 ] = 12288; 
	rom[ 2035 ] = 12288; 
	rom[ 2036 ] = 8192; 
	rom[ 2037 ] = 8192; 
	rom[ 2038 ] = 12288; 
	rom[ 2039 ] = 8192; 
	rom[ 2040 ] = 8192; 
	rom[ 2041 ] = 8192; 
	rom[ 2042 ] = 8192; 
	rom[ 2043 ] = 8192; 
	rom[ 2044 ] = 8192; 
	rom[ 2045 ] = 12288; 
	rom[ 2046 ] = 8192; 
	rom[ 2047 ] = 8192; 
	rom[ 2048 ] = 12288; 
	rom[ 2049 ] = 12288; 
	rom[ 2050 ] = 12288; 
	rom[ 2051 ] = 12288; 
	rom[ 2052 ] = 12288; 
	rom[ 2053 ] = 8192; 
	rom[ 2054 ] = 8192; 
	rom[ 2055 ] = 12288; 
	rom[ 2056 ] = 8192; 
	rom[ 2057 ] = 12288; 
	rom[ 2058 ] = 12288; 
	rom[ 2059 ] = 12288; 
	rom[ 2060 ] = 8192; 
	rom[ 2061 ] = 8192; 
	rom[ 2062 ] = 12288; 
	rom[ 2063 ] = 12288; 
	rom[ 2064 ] = 12288; 
	rom[ 2065 ] = 12288; 
	rom[ 2066 ] = 12288; 
	rom[ 2067 ] = 8192; 
	rom[ 2068 ] = 8192; 
	rom[ 2069 ] = 8192; 
	rom[ 2070 ] = 8192; 
	rom[ 2071 ] = 8192; 
	rom[ 2072 ] = 8192; 
	rom[ 2073 ] = 8192; 
	rom[ 2074 ] = 8192; 
	rom[ 2075 ] = 12288; 
	rom[ 2076 ] = 8192; 
	rom[ 2077 ] = 12288; 
	rom[ 2078 ] = 8192; 
	rom[ 2079 ] = 12288; 
	rom[ 2080 ] = 8192; 
	rom[ 2081 ] = 8192; 
	rom[ 2082 ] = 8192; 
	rom[ 2083 ] = 8192; 
	rom[ 2084 ] = 8192; 
	rom[ 2085 ] = 12288; 
	rom[ 2086 ] = 12288; 
	rom[ 2087 ] = 12288; 
	rom[ 2088 ] = 12288; 
	rom[ 2089 ] = 8192; 
	rom[ 2090 ] = 8192; 
	rom[ 2091 ] = 8192; 
	rom[ 2092 ] = 8192; 
	rom[ 2093 ] = 12288; 
	rom[ 2094 ] = 8192; 
	rom[ 2095 ] = 8192; 
	rom[ 2096 ] = 8192; 
	rom[ 2097 ] = 12288; 
	rom[ 2098 ] = 12288; 
	rom[ 2099 ] = 8192; 
	rom[ 2100 ] = 12288; 
	rom[ 2101 ] = 12288; 
	rom[ 2102 ] = 8192; 
	rom[ 2103 ] = 8192; 
	rom[ 2104 ] = 8192; 
	rom[ 2105 ] = 8192; 
	rom[ 2106 ] = 8192; 
	rom[ 2107 ] = 12288; 
	rom[ 2108 ] = 8192; 
	rom[ 2109 ] = 8192; 
	rom[ 2110 ] = 8192; 
	rom[ 2111 ] = 12288; 
	rom[ 2112 ] = 8192; 
	rom[ 2113 ] = 8192; 
	rom[ 2114 ] = 8192; 
	rom[ 2115 ] = 8192; 
	rom[ 2116 ] = 12288; 
	rom[ 2117 ] = 8192; 
	rom[ 2118 ] = 12288; 
	rom[ 2119 ] = 12288; 
	rom[ 2120 ] = 12288; 
	rom[ 2121 ] = 12288; 
	rom[ 2122 ] = 12288; 
	rom[ 2123 ] = 12288; 
	rom[ 2124 ] = 12288; 
	rom[ 2125 ] = 12288; 
	rom[ 2126 ] = 12288; 
	rom[ 2127 ] = 8192; 
	rom[ 2128 ] = 12288; 
	rom[ 2129 ] = 12288; 
	rom[ 2130 ] = 12288; 
	rom[ 2131 ] = 8192; 
	rom[ 2132 ] = 8192; 
	rom[ 2133 ] = 8192; 
	rom[ 2134 ] = 12288; 
	rom[ 2135 ] = 8192; 
	rom[ 2136 ] = 12288; 
	rom[ 2137 ] = 8192; 
	rom[ 2138 ] = 8192; 
	rom[ 2139 ] = 12288; 
	rom[ 2140 ] = 12288; 
	rom[ 2141 ] = 8192; 
	rom[ 2142 ] = 8192; 
	rom[ 2143 ] = 12288; 
	rom[ 2144 ] = 12288; 
	rom[ 2145 ] = 12288; 
	rom[ 2146 ] = 8192; 
	rom[ 2147 ] = 8192; 
	rom[ 2148 ] = 8192; 
	rom[ 2149 ] = 12288; 
	rom[ 2150 ] = 12288; 
	rom[ 2151 ] = 12288; 
	rom[ 2152 ] = 12288; 
	rom[ 2153 ] = 8192; 
	rom[ 2154 ] = 12288; 
	rom[ 2155 ] = 8192; 
	rom[ 2156 ] = 8192; 
	rom[ 2157 ] = 8192; 
	rom[ 2158 ] = 12288; 
	rom[ 2159 ] = 12288; 
	rom[ 2160 ] = 12288; 
	rom[ 2161 ] = 12288; 
	rom[ 2162 ] = 12288; 
	rom[ 2163 ] = 12288; 
	rom[ 2164 ] = 8192; 
	rom[ 2165 ] = 8192; 
	rom[ 2166 ] = 8192; 
	rom[ 2167 ] = 8192; 
	rom[ 2168 ] = 12288; 
	rom[ 2169 ] = 12288; 
	rom[ 2170 ] = 8192; 
	rom[ 2171 ] = 12288; 
	rom[ 2172 ] = 12288; 
	rom[ 2173 ] = 12288; 
	rom[ 2174 ] = 8192; 
	rom[ 2175 ] = 12288; 
	rom[ 2176 ] = 12288; 
	rom[ 2177 ] = 8192; 
	rom[ 2178 ] = 8192; 
	rom[ 2179 ] = 12288; 
	rom[ 2180 ] = 12288; 
	rom[ 2181 ] = 8192; 
	rom[ 2182 ] = 12288; 
	rom[ 2183 ] = 12288; 
	rom[ 2184 ] = 12288; 
	rom[ 2185 ] = 12288; 
	rom[ 2186 ] = 8192; 
	rom[ 2187 ] = 12288; 
	rom[ 2188 ] = 12288; 
	rom[ 2189 ] = 8192; 
	rom[ 2190 ] = 8192; 
	rom[ 2191 ] = 8192; 
	rom[ 2192 ] = 8192; 
	rom[ 2193 ] = 12288; 
	rom[ 2194 ] = 12288; 
	rom[ 2195 ] = 12288; 
	rom[ 2196 ] = 12288; 
	rom[ 2197 ] = 8192; 
	rom[ 2198 ] = 12288; 
	rom[ 2199 ] = 8192; 
	rom[ 2200 ] = 12288; 
	rom[ 2201 ] = 12288; 
	rom[ 2202 ] = 8192; 
	rom[ 2203 ] = 12288; 
	rom[ 2204 ] = 8192; 
	rom[ 2205 ] = 8192; 
	rom[ 2206 ] = 8192; 
	rom[ 2207 ] = 12288; 
	rom[ 2208 ] = 12288; 
	rom[ 2209 ] = 12288; 
	rom[ 2210 ] = 12288; 
	rom[ 2211 ] = 12288; 
	rom[ 2212 ] = 12288; 
	rom[ 2213 ] = 8192; 
	rom[ 2214 ] = 8192; 
	rom[ 2215 ] = 12288; 
	rom[ 2216 ] = 12288; 
	rom[ 2217 ] = 12288; 
	rom[ 2218 ] = 8192; 
	rom[ 2219 ] = 12288; 
	rom[ 2220 ] = 12288; 
	rom[ 2221 ] = 12288; 
	rom[ 2222 ] = 12288; 
	rom[ 2223 ] = 12288; 
	rom[ 2224 ] = 12288; 
	rom[ 2225 ] = 8192; 
	rom[ 2226 ] = 8192; 
	rom[ 2227 ] = 12288; 
	rom[ 2228 ] = 12288; 
	rom[ 2229 ] = 12288; 
	rom[ 2230 ] = 8192; 
	rom[ 2231 ] = 12288; 
	rom[ 2232 ] = 12288; 
	rom[ 2233 ] = 12288; 
	rom[ 2234 ] = 12288; 
	rom[ 2235 ] = 12288; 
	rom[ 2236 ] = 12288; 
	rom[ 2237 ] = 8192; 
	rom[ 2238 ] = 8192; 
	rom[ 2239 ] = 8192; 
	rom[ 2240 ] = 8192; 
	rom[ 2241 ] = 12288; 
	rom[ 2242 ] = 8192; 
	rom[ 2243 ] = 8192; 
	rom[ 2244 ] = 8192; 
	rom[ 2245 ] = 8192; 
	rom[ 2246 ] = 8192; 
	rom[ 2247 ] = 8192; 
	rom[ 2248 ] = 8192; 
	rom[ 2249 ] = 12288; 
	rom[ 2250 ] = 8192; 
	rom[ 2251 ] = 12288; 
	rom[ 2252 ] = 8192; 
	rom[ 2253 ] = 8192; 
	rom[ 2254 ] = 12288; 
	rom[ 2255 ] = 8192; 
	rom[ 2256 ] = 12288; 
	rom[ 2257 ] = 12288; 
	rom[ 2258 ] = 12288; 
	rom[ 2259 ] = 12288; 
	rom[ 2260 ] = 12288; 
	rom[ 2261 ] = 12288; 
	rom[ 2262 ] = 12288; 
	rom[ 2263 ] = 8192; 
	rom[ 2264 ] = 8192; 
	rom[ 2265 ] = 8192; 
	rom[ 2266 ] = 8192; 
	rom[ 2267 ] = 12288; 
	rom[ 2268 ] = 12288; 
	rom[ 2269 ] = 8192; 
	rom[ 2270 ] = 8192; 
	rom[ 2271 ] = 8192; 
	rom[ 2272 ] = 8192; 
	rom[ 2273 ] = 8192; 
	rom[ 2274 ] = 8192; 
	rom[ 2275 ] = 8192; 
	rom[ 2276 ] = 12288; 
	rom[ 2277 ] = 8192; 
	rom[ 2278 ] = 8192; 
	rom[ 2279 ] = 8192; 
	rom[ 2280 ] = 12288; 
	rom[ 2281 ] = 8192; 
	rom[ 2282 ] = 12288; 
	rom[ 2283 ] = 12288; 
	rom[ 2284 ] = 12288; 
	rom[ 2285 ] = 12288; 
	rom[ 2286 ] = 8192; 
	rom[ 2287 ] = 8192; 
	rom[ 2288 ] = 12288; 
	rom[ 2289 ] = 8192; 
	rom[ 2290 ] = 8192; 
	rom[ 2291 ] = 8192; 
	rom[ 2292 ] = 8192; 
	rom[ 2293 ] = 12288; 
	rom[ 2294 ] = 12288; 
	rom[ 2295 ] = 8192; 
	rom[ 2296 ] = 8192; 
	rom[ 2297 ] = 12288; 
	rom[ 2298 ] = 8192; 
	rom[ 2299 ] = 8192; 
	rom[ 2300 ] = 8192; 
	rom[ 2301 ] = 12288; 
	rom[ 2302 ] = 12288; 
	rom[ 2303 ] = 12288; 
	rom[ 2304 ] = 12288; 
	rom[ 2305 ] = 8192; 
	rom[ 2306 ] = 8192; 
	rom[ 2307 ] = 12288; 
	rom[ 2308 ] = 12288; 
	rom[ 2309 ] = 12288; 
	rom[ 2310 ] = 12288; 
	rom[ 2311 ] = 12288; 
	rom[ 2312 ] = 12288; 
	rom[ 2313 ] = 12288; 
	rom[ 2314 ] = 12288; 
	rom[ 2315 ] = 12288; 
	rom[ 2316 ] = 12288; 
	rom[ 2317 ] = 8192; 
	rom[ 2318 ] = 8192; 
	rom[ 2319 ] = 8192; 
	rom[ 2320 ] = 8192; 
	rom[ 2321 ] = 8192; 
	rom[ 2322 ] = 8192; 
	rom[ 2323 ] = 8192; 
	rom[ 2324 ] = 12288; 
	rom[ 2325 ] = 8192; 
	rom[ 2326 ] = 8192; 
	rom[ 2327 ] = 12288; 
	rom[ 2328 ] = 12288; 
	rom[ 2329 ] = 8192; 
	rom[ 2330 ] = 12288; 
	rom[ 2331 ] = 8192; 
	rom[ 2332 ] = 8192; 
	rom[ 2333 ] = 12288; 
	rom[ 2334 ] = 12288; 
	rom[ 2335 ] = 12288; 
	rom[ 2336 ] = 12288; 
	rom[ 2337 ] = 8192; 
	rom[ 2338 ] = 8192; 
	rom[ 2339 ] = 8192; 
	rom[ 2340 ] = 12288; 
	rom[ 2341 ] = 8192; 
	rom[ 2342 ] = 12288; 
	rom[ 2343 ] = 12288; 
	rom[ 2344 ] = 12288; 
	rom[ 2345 ] = 12288; 
	rom[ 2346 ] = 8192; 
	rom[ 2347 ] = 8192; 
	rom[ 2348 ] = 8192; 
	rom[ 2349 ] = 8192; 
	rom[ 2350 ] = 8192; 
	rom[ 2351 ] = 8192; 
	rom[ 2352 ] = 12288; 
	rom[ 2353 ] = 12288; 
	rom[ 2354 ] = 8192; 
	rom[ 2355 ] = 12288; 
	rom[ 2356 ] = 8192; 
	rom[ 2357 ] = 8192; 
	rom[ 2358 ] = 8192; 
	rom[ 2359 ] = 8192; 
	rom[ 2360 ] = 8192; 
	rom[ 2361 ] = 8192; 
	rom[ 2362 ] = 12288; 
	rom[ 2363 ] = 12288; 
	rom[ 2364 ] = 12288; 
	rom[ 2365 ] = 8192; 
	rom[ 2366 ] = 12288; 
	rom[ 2367 ] = 12288; 
	rom[ 2368 ] = 8192; 
	rom[ 2369 ] = 8192; 
	rom[ 2370 ] = 8192; 
	rom[ 2371 ] = 8192; 
	rom[ 2372 ] = 8192; 
	rom[ 2373 ] = 12288; 
	rom[ 2374 ] = 8192; 
	rom[ 2375 ] = 12288; 
	rom[ 2376 ] = 8192; 
	rom[ 2377 ] = 8192; 
	rom[ 2378 ] = 8192; 
	rom[ 2379 ] = 12288; 
	rom[ 2380 ] = 12288; 
	rom[ 2381 ] = 8192; 
	rom[ 2382 ] = 8192; 
	rom[ 2383 ] = 8192; 
	rom[ 2384 ] = 8192; 
	rom[ 2385 ] = 8192; 
	rom[ 2386 ] = 8192; 
	rom[ 2387 ] = 8192; 
	rom[ 2388 ] = 8192; 
	rom[ 2389 ] = 12288; 
	rom[ 2390 ] = 12288; 
	rom[ 2391 ] = 8192; 
	rom[ 2392 ] = 8192; 
	rom[ 2393 ] = 8192; 
	rom[ 2394 ] = 12288; 
	rom[ 2395 ] = 8192; 
	rom[ 2396 ] = 12288; 
	rom[ 2397 ] = 12288; 
	rom[ 2398 ] = 12288; 
	rom[ 2399 ] = 12288; 
	rom[ 2400 ] = 8192; 
	rom[ 2401 ] = 8192; 
	rom[ 2402 ] = 8192; 
	rom[ 2403 ] = 12288; 
	rom[ 2404 ] = 8192; 
	rom[ 2405 ] = 8192; 
	rom[ 2406 ] = 12288; 
	rom[ 2407 ] = 12288; 
	rom[ 2408 ] = 12288; 
	rom[ 2409 ] = 12288; 
	rom[ 2410 ] = 12288; 
	rom[ 2411 ] = 8192; 
	rom[ 2412 ] = 8192; 
	rom[ 2413 ] = 12288; 
	rom[ 2414 ] = 12288; 
	rom[ 2415 ] = 12288; 
	rom[ 2416 ] = 8192; 
	rom[ 2417 ] = 12288; 
	rom[ 2418 ] = 12288; 
	rom[ 2419 ] = 8192; 
	rom[ 2420 ] = 8192; 
	rom[ 2421 ] = 8192; 
	rom[ 2422 ] = 12288; 
	rom[ 2423 ] = 12288; 
	rom[ 2424 ] = 12288; 
	rom[ 2425 ] = 8192; 
	rom[ 2426 ] = 12288; 
	rom[ 2427 ] = 8192; 
	rom[ 2428 ] = 8192; 
	rom[ 2429 ] = 8192; 
	rom[ 2430 ] = 12288; 
	rom[ 2431 ] = 12288; 
	rom[ 2432 ] = 12288; 
	rom[ 2433 ] = 8192; 
	rom[ 2434 ] = 8192; 
	rom[ 2435 ] = 8192; 
	rom[ 2436 ] = 8192; 
	rom[ 2437 ] = 8192; 
	rom[ 2438 ] = 8192; 
	rom[ 2439 ] = 8192; 
	rom[ 2440 ] = 12288; 
	rom[ 2441 ] = 8192; 
	rom[ 2442 ] = 12288; 
	rom[ 2443 ] = 8192; 
	rom[ 2444 ] = 8192; 
	rom[ 2445 ] = 8192; 
	rom[ 2446 ] = 12288; 
	rom[ 2447 ] = 12288; 
	rom[ 2448 ] = 8192; 
	rom[ 2449 ] = 8192; 
	rom[ 2450 ] = 12288; 
	rom[ 2451 ] = 12288; 
	rom[ 2452 ] = 8192; 
	rom[ 2453 ] = 8192; 
	rom[ 2454 ] = 8192; 
	rom[ 2455 ] = 12288; 
	rom[ 2456 ] = 8192; 
	rom[ 2457 ] = 8192; 
	rom[ 2458 ] = 12288; 
	rom[ 2459 ] = 12288; 
	rom[ 2460 ] = 8192; 
	rom[ 2461 ] = 12288; 
	rom[ 2462 ] = 8192; 
	rom[ 2463 ] = 8192; 
	rom[ 2464 ] = 12288; 
	rom[ 2465 ] = 12288; 
	rom[ 2466 ] = 12288; 
	rom[ 2467 ] = 12288; 
	rom[ 2468 ] = 12288; 
	rom[ 2469 ] = 12288; 
	rom[ 2470 ] = 12288; 
	rom[ 2471 ] = 12288; 
	rom[ 2472 ] = 12288; 
	rom[ 2473 ] = 12288; 
	rom[ 2474 ] = 12288; 
	rom[ 2475 ] = 8192; 
	rom[ 2476 ] = 8192; 
	rom[ 2477 ] = 8192; 
	rom[ 2478 ] = 12288; 
	rom[ 2479 ] = 8192; 
	rom[ 2480 ] = 12288; 
	rom[ 2481 ] = 8192; 
	rom[ 2482 ] = 8192; 
	rom[ 2483 ] = 8192; 
	rom[ 2484 ] = 12288; 
	rom[ 2485 ] = 8192; 
	rom[ 2486 ] = 12288; 
	rom[ 2487 ] = 12288; 
	rom[ 2488 ] = 12288; 
	rom[ 2489 ] = 12288; 
	rom[ 2490 ] = 8192; 
	rom[ 2491 ] = 8192; 
	rom[ 2492 ] = 8192; 
	rom[ 2493 ] = 8192; 
	rom[ 2494 ] = 8192; 
	rom[ 2495 ] = 12288; 
	rom[ 2496 ] = 8192; 
	rom[ 2497 ] = 12288; 
	rom[ 2498 ] = 12288; 
	rom[ 2499 ] = 8192; 
	rom[ 2500 ] = 12288; 
	rom[ 2501 ] = 8192; 
	rom[ 2502 ] = 12288; 
	rom[ 2503 ] = 12288; 
	rom[ 2504 ] = 8192; 
	rom[ 2505 ] = 8192; 
	rom[ 2506 ] = 8192; 
	rom[ 2507 ] = 8192; 
	rom[ 2508 ] = 8192; 
	rom[ 2509 ] = 12288; 
	rom[ 2510 ] = 8192; 
	rom[ 2511 ] = 8192; 
	rom[ 2512 ] = 12288; 
	rom[ 2513 ] = 8192; 
	rom[ 2514 ] = 12288; 
	rom[ 2515 ] = 8192; 
	rom[ 2516 ] = 8192; 
	rom[ 2517 ] = 12288; 
	rom[ 2518 ] = 12288; 
	rom[ 2519 ] = 12288; 
	rom[ 2520 ] = 12288; 
	rom[ 2521 ] = 12288; 
	rom[ 2522 ] = 12288; 
	rom[ 2523 ] = 12288; 
	rom[ 2524 ] = 12288; 
	rom[ 2525 ] = 12288; 
	rom[ 2526 ] = 12288; 
	rom[ 2527 ] = 8192; 
	rom[ 2528 ] = 8192; 
	rom[ 2529 ] = 12288; 
	rom[ 2530 ] = 8192; 
	rom[ 2531 ] = 8192; 
	rom[ 2532 ] = 8192; 
	rom[ 2533 ] = 12288; 
	rom[ 2534 ] = 12288; 
	rom[ 2535 ] = 8192; 
	rom[ 2536 ] = 8192; 
	rom[ 2537 ] = 8192; 
	rom[ 2538 ] = 12288; 
	rom[ 2539 ] = 8192; 
	rom[ 2540 ] = 8192; 
	rom[ 2541 ] = 12288; 
	rom[ 2542 ] = 8192; 
	rom[ 2543 ] = 8192; 
	rom[ 2544 ] = 8192; 
	rom[ 2545 ] = 12288; 
	rom[ 2546 ] = 12288; 
	rom[ 2547 ] = 12288; 
	rom[ 2548 ] = 12288; 
	rom[ 2549 ] = 12288; 
	rom[ 2550 ] = 8192; 
	rom[ 2551 ] = 12288; 
	rom[ 2552 ] = 12288; 
	rom[ 2553 ] = 8192; 
	rom[ 2554 ] = 12288; 
	rom[ 2555 ] = 8192; 
	rom[ 2556 ] = 12288; 
	rom[ 2557 ] = 8192; 
	rom[ 2558 ] = 8192; 
	rom[ 2559 ] = 8192; 
	rom[ 2560 ] = 12288; 
	rom[ 2561 ] = 8192; 
	rom[ 2562 ] = 8192; 
	rom[ 2563 ] = 12288; 
	rom[ 2564 ] = 12288; 
	rom[ 2565 ] = 12288; 
	rom[ 2566 ] = 12288; 
	rom[ 2567 ] = 12288; 
	rom[ 2568 ] = 8192; 
	rom[ 2569 ] = 8192; 
	rom[ 2570 ] = 12288; 
	rom[ 2571 ] = 12288; 
	rom[ 2572 ] = 8192; 
	rom[ 2573 ] = 8192; 
	rom[ 2574 ] = 12288; 
	rom[ 2575 ] = 12288; 
	rom[ 2576 ] = 12288; 
	rom[ 2577 ] = 12288; 
	rom[ 2578 ] = 12288; 
	rom[ 2579 ] = 12288; 
	rom[ 2580 ] = 8192; 
	rom[ 2581 ] = 8192; 
	rom[ 2582 ] = 8192; 
	rom[ 2583 ] = 8192; 
	rom[ 2584 ] = 8192; 
	rom[ 2585 ] = 8192; 
	rom[ 2586 ] = 8192; 
	rom[ 2587 ] = 8192; 
	rom[ 2588 ] = 12288; 
	rom[ 2589 ] = 8192; 
	rom[ 2590 ] = 8192; 
	rom[ 2591 ] = 8192; 
	rom[ 2592 ] = 8192; 
	rom[ 2593 ] = 12288; 
	rom[ 2594 ] = 12288; 
	rom[ 2595 ] = 8192; 
	rom[ 2596 ] = 12288; 
	rom[ 2597 ] = 8192; 
	rom[ 2598 ] = 8192; 
	rom[ 2599 ] = 12288; 
	rom[ 2600 ] = 12288; 
	rom[ 2601 ] = 12288; 
	rom[ 2602 ] = 12288; 
	rom[ 2603 ] = 8192; 
	rom[ 2604 ] = 8192; 
	rom[ 2605 ] = 8192; 
	rom[ 2606 ] = 12288; 
	rom[ 2607 ] = 12288; 
	rom[ 2608 ] = 8192; 
	rom[ 2609 ] = 12288; 
	rom[ 2610 ] = 12288; 
	rom[ 2611 ] = 8192; 
	rom[ 2612 ] = 8192; 
	rom[ 2613 ] = 8192; 
	rom[ 2614 ] = 8192; 
	rom[ 2615 ] = 12288; 
	rom[ 2616 ] = 8192; 
	rom[ 2617 ] = 12288; 
	rom[ 2618 ] = 12288; 
	rom[ 2619 ] = 12288; 
	rom[ 2620 ] = 12288; 
	rom[ 2621 ] = 12288; 
	rom[ 2622 ] = 8192; 
	rom[ 2623 ] = 8192; 
	rom[ 2624 ] = 8192; 
	rom[ 2625 ] = 12288; 
	rom[ 2626 ] = 8192; 
	rom[ 2627 ] = 8192; 
	rom[ 2628 ] = 8192; 
	rom[ 2629 ] = 12288; 
	rom[ 2630 ] = 12288; 
	rom[ 2631 ] = 12288; 
	rom[ 2632 ] = 8192; 
	rom[ 2633 ] = 8192; 
	rom[ 2634 ] = 12288; 
	rom[ 2635 ] = 8192; 
	rom[ 2636 ] = 8192; 
	rom[ 2637 ] = 8192; 
	rom[ 2638 ] = 12288; 
	rom[ 2639 ] = 8192; 
	rom[ 2640 ] = 12288; 
	rom[ 2641 ] = 8192; 
	rom[ 2642 ] = 8192; 
	rom[ 2643 ] = 8192; 
	rom[ 2644 ] = 12288; 
	rom[ 2645 ] = 8192; 
	rom[ 2646 ] = 8192; 
	rom[ 2647 ] = 8192; 
	rom[ 2648 ] = 8192; 
	rom[ 2649 ] = 8192; 
	rom[ 2650 ] = 8192; 
	rom[ 2651 ] = 12288; 
	rom[ 2652 ] = 12288; 
	rom[ 2653 ] = 8192; 
	rom[ 2654 ] = 12288; 
	rom[ 2655 ] = 12288; 
	rom[ 2656 ] = 8192; 
	rom[ 2657 ] = 12288; 
	rom[ 2658 ] = 12288; 
	rom[ 2659 ] = 12288; 
	rom[ 2660 ] = 12288; 
	rom[ 2661 ] = 12288; 
	rom[ 2662 ] = 12288; 
	rom[ 2663 ] = 12288; 
	rom[ 2664 ] = 12288; 
	rom[ 2665 ] = 8192; 
	rom[ 2666 ] = 8192; 
	rom[ 2667 ] = 12288; 
	rom[ 2668 ] = 12288; 
	rom[ 2669 ] = 12288; 
	rom[ 2670 ] = 8192; 
	rom[ 2671 ] = 8192; 
	rom[ 2672 ] = 12288; 
	rom[ 2673 ] = 12288; 
	rom[ 2674 ] = 8192; 
	rom[ 2675 ] = 8192; 
	rom[ 2676 ] = 8192; 
	rom[ 2677 ] = 12288; 
	rom[ 2678 ] = 12288; 
	rom[ 2679 ] = 8192; 
	rom[ 2680 ] = 12288; 
	rom[ 2681 ] = 8192; 
	rom[ 2682 ] = 8192; 
	rom[ 2683 ] = 12288; 
	rom[ 2684 ] = 12288; 
	rom[ 2685 ] = 8192; 
	rom[ 2686 ] = 8192; 
	rom[ 2687 ] = 12288; 
	rom[ 2688 ] = 12288; 
	rom[ 2689 ] = 8192; 
	rom[ 2690 ] = 12288; 
	rom[ 2691 ] = 8192; 
	rom[ 2692 ] = 12288; 
	rom[ 2693 ] = 8192; 
	rom[ 2694 ] = 8192; 
	rom[ 2695 ] = 12288; 
	rom[ 2696 ] = 12288; 
	rom[ 2697 ] = 12288; 
	rom[ 2698 ] = 12288; 
	rom[ 2699 ] = 12288; 
	rom[ 2700 ] = 12288; 
	rom[ 2701 ] = 12288; 
	rom[ 2702 ] = 12288; 
	rom[ 2703 ] = 8192; 
	rom[ 2704 ] = 8192; 
	rom[ 2705 ] = 8192; 
	rom[ 2706 ] = 8192; 
	rom[ 2707 ] = 8192; 
	rom[ 2708 ] = 12288; 
	rom[ 2709 ] = 12288; 
	rom[ 2710 ] = 12288; 
	rom[ 2711 ] = 8192; 
	rom[ 2712 ] = 8192; 
	rom[ 2713 ] = 12288; 
	rom[ 2714 ] = 12288; 
	rom[ 2715 ] = 8192; 
	rom[ 2716 ] = 8192; 
	rom[ 2717 ] = 12288; 
	rom[ 2718 ] = 8192; 
	rom[ 2719 ] = 8192; 
	rom[ 2720 ] = 8192; 
	rom[ 2721 ] = 12288; 
	rom[ 2722 ] = 8192; 
	rom[ 2723 ] = 8192; 
	rom[ 2724 ] = 12288; 
	rom[ 2725 ] = 12288; 
	rom[ 2726 ] = 12288; 
	rom[ 2727 ] = 12288; 
	rom[ 2728 ] = 8192; 
	rom[ 2729 ] = 8192; 
	rom[ 2730 ] = 12288; 
	rom[ 2731 ] = 8192; 
	rom[ 2732 ] = 8192; 
	rom[ 2733 ] = 12288; 
	rom[ 2734 ] = 12288; 
	rom[ 2735 ] = 12288; 
	rom[ 2736 ] = 8192; 
	rom[ 2737 ] = 12288; 
	rom[ 2738 ] = 8192; 
	rom[ 2739 ] = 12288; 
	rom[ 2740 ] = 12288; 
	rom[ 2741 ] = 12288; 
	rom[ 2742 ] = 12288; 
	rom[ 2743 ] = 12288; 
	rom[ 2744 ] = 8192; 
	rom[ 2745 ] = 8192; 
	rom[ 2746 ] = 12288; 
	rom[ 2747 ] = 8192; 
	rom[ 2748 ] = 8192; 
	rom[ 2749 ] = 8192; 
	rom[ 2750 ] = 8192; 
	rom[ 2751 ] = 8192; 
	rom[ 2752 ] = 12288; 
	rom[ 2753 ] = 12288; 
	rom[ 2754 ] = 12288; 
	rom[ 2755 ] = 8192; 
	rom[ 2756 ] = 8192; 
	rom[ 2757 ] = 8192; 
	rom[ 2758 ] = 12288; 
	rom[ 2759 ] = 8192; 
	rom[ 2760 ] = 12288; 
	rom[ 2761 ] = 8192; 
	rom[ 2762 ] = 8192; 
	rom[ 2763 ] = 8192; 
	rom[ 2764 ] = 12288; 
	rom[ 2765 ] = 12288; 
	rom[ 2766 ] = 12288; 
	rom[ 2767 ] = 12288; 
	rom[ 2768 ] = 12288; 
	rom[ 2769 ] = 8192; 
	rom[ 2770 ] = 8192; 
	rom[ 2771 ] = 8192; 
	rom[ 2772 ] = 12288; 
	rom[ 2773 ] = 8192; 
	rom[ 2774 ] = 8192; 
	rom[ 2775 ] = 8192; 
	rom[ 2776 ] = 8192; 
	rom[ 2777 ] = 8192; 
	rom[ 2778 ] = 8192; 
	rom[ 2779 ] = 8192; 
	rom[ 2780 ] = 12288; 
	rom[ 2781 ] = 12288; 
	rom[ 2782 ] = 12288; 
	rom[ 2783 ] = 12288; 
	rom[ 2784 ] = 8192; 
	rom[ 2785 ] = 12288; 
	rom[ 2786 ] = 8192; 
	rom[ 2787 ] = 12288; 
	rom[ 2788 ] = 12288; 
	rom[ 2789 ] = 8192; 
	rom[ 2790 ] = 8192; 
	rom[ 2791 ] = 8192; 
	rom[ 2792 ] = 8192; 
	rom[ 2793 ] = 8192; 
	rom[ 2794 ] = 8192; 
	rom[ 2795 ] = 8192; 
	rom[ 2796 ] = 12288; 
	rom[ 2797 ] = 8192; 
	rom[ 2798 ] = 8192; 
	rom[ 2799 ] = 8192; 
	rom[ 2800 ] = 8192; 
	rom[ 2801 ] = 8192; 
	rom[ 2802 ] = 12288; 
	rom[ 2803 ] = 12288; 
	rom[ 2804 ] = 12288; 
	rom[ 2805 ] = 12288; 
	rom[ 2806 ] = 12288; 
	rom[ 2807 ] = 12288; 
	rom[ 2808 ] = 12288; 
	rom[ 2809 ] = 12288; 
	rom[ 2810 ] = 12288; 
	rom[ 2811 ] = 12288; 
	rom[ 2812 ] = 12288; 
	rom[ 2813 ] = 8192; 
	rom[ 2814 ] = 8192; 
	rom[ 2815 ] = 8192; 
	rom[ 2816 ] = 8192; 
	rom[ 2817 ] = 8192; 
	rom[ 2818 ] = 8192; 
	rom[ 2819 ] = 12288; 
	rom[ 2820 ] = 8192; 
	rom[ 2821 ] = 12288; 
	rom[ 2822 ] = 12288; 
	rom[ 2823 ] = 12288; 
	rom[ 2824 ] = 12288; 
	rom[ 2825 ] = 12288; 
	rom[ 2826 ] = 8192; 
	rom[ 2827 ] = 12288; 
	rom[ 2828 ] = 12288; 
	rom[ 2829 ] = 12288; 
	rom[ 2830 ] = 12288; 
	rom[ 2831 ] = 8192; 
	rom[ 2832 ] = 8192; 
	rom[ 2833 ] = 12288; 
	rom[ 2834 ] = 12288; 
	rom[ 2835 ] = 12288; 
	rom[ 2836 ] = 12288; 
	rom[ 2837 ] = 8192; 
	rom[ 2838 ] = 8192; 
	rom[ 2839 ] = 12288; 
	rom[ 2840 ] = 12288; 
	rom[ 2841 ] = 12288; 
	rom[ 2842 ] = 12288; 
	rom[ 2843 ] = 12288; 
	rom[ 2844 ] = 12288; 
	rom[ 2845 ] = 12288; 
	rom[ 2846 ] = 8192; 
	rom[ 2847 ] = 12288; 
	rom[ 2848 ] = 12288; 
	rom[ 2849 ] = 12288; 
	rom[ 2850 ] = 12288; 
	rom[ 2851 ] = 8192; 
	rom[ 2852 ] = 8192; 
	rom[ 2853 ] = 12288; 
	rom[ 2854 ] = 12288; 
	rom[ 2855 ] = 8192; 
	rom[ 2856 ] = 8192; 
	rom[ 2857 ] = 8192; 
	rom[ 2858 ] = 8192; 
	rom[ 2859 ] = 8192; 
	rom[ 2860 ] = 8192; 
	rom[ 2861 ] = 8192; 
	rom[ 2862 ] = 8192; 
	rom[ 2863 ] = 8192; 
	rom[ 2864 ] = 8192; 
	rom[ 2865 ] = 12288; 
	rom[ 2866 ] = 8192; 
	rom[ 2867 ] = 8192; 
	rom[ 2868 ] = 12288; 
	rom[ 2869 ] = 12288; 
	rom[ 2870 ] = 12288; 
	rom[ 2871 ] = 8192; 
	rom[ 2872 ] = 12288; 
	rom[ 2873 ] = 8192; 
	rom[ 2874 ] = 12288; 
	rom[ 2875 ] = 8192; 
	rom[ 2876 ] = 8192; 
	rom[ 2877 ] = 8192; 
	rom[ 2878 ] = 8192; 
	rom[ 2879 ] = 8192; 
	rom[ 2880 ] = 8192; 
	rom[ 2881 ] = 8192; 
	rom[ 2882 ] = 8192; 
	rom[ 2883 ] = 8192; 
	rom[ 2884 ] = 12288; 
	rom[ 2885 ] = 12288; 
	rom[ 2886 ] = 12288; 
	rom[ 2887 ] = 12288; 
	rom[ 2888 ] = 12288; 
	rom[ 2889 ] = 12288; 
	rom[ 2890 ] = 8192; 
	rom[ 2891 ] = 12288; 
	rom[ 2892 ] = 12288; 
	rom[ 2893 ] = 12288; 
	rom[ 2894 ] = 8192; 
	rom[ 2895 ] = 8192; 
	rom[ 2896 ] = 8192; 
	rom[ 2897 ] = 8192; 
	rom[ 2898 ] = 8192; 
	rom[ 2899 ] = 8192; 
	rom[ 2900 ] = 12288; 
	rom[ 2901 ] = 8192; 
	rom[ 2902 ] = 12288; 
	rom[ 2903 ] = 8192; 
	rom[ 2904 ] = 12288; 
	rom[ 2905 ] = 12288; 
	rom[ 2906 ] = 12288; 
	rom[ 2907 ] = 12288; 
	rom[ 2908 ] = 12288; 
	rom[ 2909 ] = 12288; 
	rom[ 2910 ] = 12288; 
	rom[ 2911 ] = 8192; 
	rom[ 2912 ] = 8192; 
	end
endmodule
module rect2_wieght_rom(
	input 				clk,
	input		[11:0]	addr,
	output reg	[14:0]	q    // x y w h 5bit*4
	);
	reg					[14:0]	rom [4095:0];
	always @(posedge clk) q <= rom[addr];
	initial begin
		rom[ 0    ] = 0; 
		rom[ 1    ] = 0; 
		rom[ 2    ] = 0; 
		rom[ 3    ] = 0; 
		rom[ 4    ] = 0; 
		rom[ 5    ] = 0; 
		rom[ 6    ] = 0; 
		rom[ 7    ] = 0; 
		rom[ 8    ] = 0; 
		rom[ 9    ] = 0; 
		rom[ 10   ] = 0; 
		rom[ 11   ] = 0; 
		rom[ 12   ] = 0; 
		rom[ 13   ] = 0; 
		rom[ 14   ] = 0; 
		rom[ 15   ] = 0; 
		rom[ 16   ] = 0; 
		rom[ 17   ] = 0; 
		rom[ 18   ] = 0; 
		rom[ 19   ] = 0; 
		rom[ 20   ] = 0; 
		rom[ 21   ] = 0; 
		rom[ 22   ] = 0; 
		rom[ 23   ] = 0; 
		rom[ 24   ] = 0; 
		rom[ 25   ] = 0; 
		rom[ 26   ] = 0; 
		rom[ 27   ] = 0; 
		rom[ 28   ] = 0; 
		rom[ 29   ] = 0; 
		rom[ 30   ] = 0; 
		rom[ 31   ] = 0; 
		rom[ 32   ] = 0; 
		rom[ 33   ] = 0; 
		rom[ 34   ] = 0; 
		rom[ 35   ] = 8192; 
		rom[ 36   ] = 0; 
		rom[ 37   ] = 0; 
		rom[ 38   ] = 0; 
		rom[ 39   ] = 0; 
		rom[ 40   ] = 0; 
		rom[ 41   ] = 0; 
		rom[ 42   ] = 0; 
		rom[ 43   ] = 0; 
		rom[ 44   ] = 0; 
		rom[ 45   ] = 0; 
		rom[ 46   ] = 0; 
		rom[ 47   ] = 0; 
		rom[ 48   ] = 8192; 
		rom[ 49   ] = 0; 
		rom[ 50   ] = 0; 
		rom[ 51   ] = 0; 
		rom[ 52   ] = 0; 
		rom[ 53   ] = 0; 
		rom[ 54   ] = 0; 
		rom[ 55   ] = 0; 
		rom[ 56   ] = 8192; 
		rom[ 57   ] = 0; 
		rom[ 58   ] = 0; 
		rom[ 59   ] = 0; 
		rom[ 60   ] = 0; 
		rom[ 61   ] = 0; 
		rom[ 62   ] = 8192; 
		rom[ 63   ] = 0; 
		rom[ 64   ] = 0; 
		rom[ 65   ] = 0; 
		rom[ 66   ] = 0; 
		rom[ 67   ] = 0; 
		rom[ 68   ] = 0; 
		rom[ 69   ] = 0; 
		rom[ 70   ] = 8192; 
		rom[ 71   ] = 0; 
		rom[ 72   ] = 0; 
		rom[ 73   ] = 0; 
		rom[ 74   ] = 0; 
		rom[ 75   ] = 8192; 
		rom[ 76   ] = 8192; 
		rom[ 77   ] = 0; 
		rom[ 78   ] = 0; 
		rom[ 79   ] = 0; 
		rom[ 80   ] = 0; 
		rom[ 81   ] = 0; 
		rom[ 82   ] = 0; 
		rom[ 83   ] = 0; 
		rom[ 84   ] = 0; 
		rom[ 85   ] = 0; 
		rom[ 86   ] = 0; 
		rom[ 87   ] = 0; 
		rom[ 88   ] = 0; 
		rom[ 89   ] = 0; 
		rom[ 90   ] = 0; 
		rom[ 91   ] = 0; 
		rom[ 92   ] = 0; 
		rom[ 93   ] = 0; 
		rom[ 94   ] = 0; 
		rom[ 95   ] = 0; 
		rom[ 96   ] = 0; 
		rom[ 97   ] = 0; 
		rom[ 98   ] = 0; 
		rom[ 99   ] = 0; 
		rom[ 100  ] = 0; 
		rom[ 101  ] = 0; 
		rom[ 102  ] = 0; 
		rom[ 103  ] = 0; 
		rom[ 104  ] = 0; 
		rom[ 105  ] = 8192; 
		rom[ 106  ] = 0; 
		rom[ 107  ] = 0; 
		rom[ 108  ] = 0; 
		rom[ 109  ] = 8192; 
		rom[ 110  ] = 8192; 
		rom[ 111  ] = 0; 
		rom[ 112  ] = 0; 
		rom[ 113  ] = 0; 
		rom[ 114  ] = 0; 
		rom[ 115  ] = 0; 
		rom[ 116  ] = 0; 
		rom[ 117  ] = 0; 
		rom[ 118  ] = 8192; 
		rom[ 119  ] = 0; 
		rom[ 120  ] = 8192; 
		rom[ 121  ] = 8192; 
		rom[ 122  ] = 8192; 
		rom[ 123  ] = 0; 
		rom[ 124  ] = 0; 
		rom[ 125  ] = 0; 
		rom[ 126  ] = 0; 
		rom[ 127  ] = 0; 
		rom[ 128  ] = 0; 
		rom[ 129  ] = 0; 
		rom[ 130  ] = 0; 
		rom[ 131  ] = 0; 
		rom[ 132  ] = 0; 
		rom[ 133  ] = 0; 
		rom[ 134  ] = 0; 
		rom[ 135  ] = 0; 
		rom[ 136  ] = 0; 
		rom[ 137  ] = 0; 
		rom[ 138  ] = 0; 
		rom[ 139  ] = 0; 
		rom[ 140  ] = 0; 
		rom[ 141  ] = 0; 
		rom[ 142  ] = 0; 
		rom[ 143  ] = 0; 
		rom[ 144  ] = 0; 
		rom[ 145  ] = 0; 
		rom[ 146  ] = 0; 
		rom[ 147  ] = 0; 
		rom[ 148  ] = 0; 
		rom[ 149  ] = 0; 
		rom[ 150  ] = 0; 
		rom[ 151  ] = 0; 
		rom[ 152  ] = 8192; 
		rom[ 153  ] = 0; 
		rom[ 154  ] = 0; 
		rom[ 155  ] = 0; 
		rom[ 156  ] = 0; 
		rom[ 157  ] = 0; 
		rom[ 158  ] = 0; 
		rom[ 159  ] = 0; 
		rom[ 160  ] = 8192; 
		rom[ 161  ] = 0; 
		rom[ 162  ] = 0; 
		rom[ 163  ] = 0; 
		rom[ 164  ] = 8192; 
		rom[ 165  ] = 0; 
		rom[ 166  ] = 0; 
		rom[ 167  ] = 0; 
		rom[ 168  ] = 0; 
		rom[ 169  ] = 0; 
		rom[ 170  ] = 0; 
		rom[ 171  ] = 0; 
		rom[ 172  ] = 0; 
		rom[ 173  ] = 0; 
		rom[ 174  ] = 0; 
		rom[ 175  ] = 0; 
		rom[ 176  ] = 8192; 
		rom[ 177  ] = 8192; 
		rom[ 178  ] = 0; 
		rom[ 179  ] = 0; 
		rom[ 180  ] = 0; 
		rom[ 181  ] = 0; 
		rom[ 182  ] = 0; 
		rom[ 183  ] = 0; 
		rom[ 184  ] = 0; 
		rom[ 185  ] = 0; 
		rom[ 186  ] = 0; 
		rom[ 187  ] = 8192; 
		rom[ 188  ] = 0; 
		rom[ 189  ] = 0; 
		rom[ 190  ] = 0; 
		rom[ 191  ] = 0; 
		rom[ 192  ] = 0; 
		rom[ 193  ] = 0; 
		rom[ 194  ] = 0; 
		rom[ 195  ] = 0; 
		rom[ 196  ] = 0; 
		rom[ 197  ] = 0; 
		rom[ 198  ] = 0; 
		rom[ 199  ] = 0; 
		rom[ 200  ] = 0; 
		rom[ 201  ] = 0; 
		rom[ 202  ] = 8192; 
		rom[ 203  ] = 0; 
		rom[ 204  ] = 0; 
		rom[ 205  ] = 0; 
		rom[ 206  ] = 8192; 
		rom[ 207  ] = 8192; 
		rom[ 208  ] = 0; 
		rom[ 209  ] = 0; 
		rom[ 210  ] = 0; 
		rom[ 211  ] = 0; 
		rom[ 212  ] = 0; 
		rom[ 213  ] = 0; 
		rom[ 214  ] = 0; 
		rom[ 215  ] = 8192; 
		rom[ 216  ] = 0; 
		rom[ 217  ] = 8192; 
		rom[ 218  ] = 0; 
		rom[ 219  ] = 0; 
		rom[ 220  ] = 0; 
		rom[ 221  ] = 0; 
		rom[ 222  ] = 0; 
		rom[ 223  ] = 8192; 
		rom[ 224  ] = 8192; 
		rom[ 225  ] = 0; 
		rom[ 226  ] = 0; 
		rom[ 227  ] = 0; 
		rom[ 228  ] = 0; 
		rom[ 229  ] = 0; 
		rom[ 230  ] = 8192; 
		rom[ 231  ] = 0; 
		rom[ 232  ] = 0; 
		rom[ 233  ] = 0; 
		rom[ 234  ] = 8192; 
		rom[ 235  ] = 8192; 
		rom[ 236  ] = 0; 
		rom[ 237  ] = 0; 
		rom[ 238  ] = 0; 
		rom[ 239  ] = 0; 
		rom[ 240  ] = 0; 
		rom[ 241  ] = 8192; 
		rom[ 242  ] = 8192; 
		rom[ 243  ] = 0; 
		rom[ 244  ] = 0; 
		rom[ 245  ] = 0; 
		rom[ 246  ] = 0; 
		rom[ 247  ] = 0; 
		rom[ 248  ] = 8192; 
		rom[ 249  ] = 8192; 
		rom[ 250  ] = 0; 
		rom[ 251  ] = 0; 
		rom[ 252  ] = 0; 
		rom[ 253  ] = 0; 
		rom[ 254  ] = 0; 
		rom[ 255  ] = 8192; 
		rom[ 256  ] = 0; 
		rom[ 257  ] = 0; 
		rom[ 258  ] = 0; 
		rom[ 259  ] = 0; 
		rom[ 260  ] = 0; 
		rom[ 261  ] = 8192; 
		rom[ 262  ] = 0; 
		rom[ 263  ] = 0; 
		rom[ 264  ] = 0; 
		rom[ 265  ] = 0; 
		rom[ 266  ] = 0; 
		rom[ 267  ] = 0; 
		rom[ 268  ] = 0; 
		rom[ 269  ] = 0; 
		rom[ 270  ] = 0; 
		rom[ 271  ] = 0; 
		rom[ 272  ] = 0; 
		rom[ 273  ] = 0; 
		rom[ 274  ] = 0; 
		rom[ 275  ] = 0; 
		rom[ 276  ] = 0; 
		rom[ 277  ] = 0; 
		rom[ 278  ] = 0; 
		rom[ 279  ] = 0; 
		rom[ 280  ] = 0; 
		rom[ 281  ] = 0; 
		rom[ 282  ] = 0; 
		rom[ 283  ] = 0; 
		rom[ 284  ] = 0; 
		rom[ 285  ] = 0; 
		rom[ 286  ] = 0; 
		rom[ 287  ] = 0; 
		rom[ 288  ] = 8192; 
		rom[ 289  ] = 0; 
		rom[ 290  ] = 0; 
		rom[ 291  ] = 8192; 
		rom[ 292  ] = 0; 
		rom[ 293  ] = 0; 
		rom[ 294  ] = 0; 
		rom[ 295  ] = 0; 
		rom[ 296  ] = 0; 
		rom[ 297  ] = 0; 
		rom[ 298  ] = 0; 
		rom[ 299  ] = 0; 
		rom[ 300  ] = 0; 
		rom[ 301  ] = 0; 
		rom[ 302  ] = 0; 
		rom[ 303  ] = 0; 
		rom[ 304  ] = 0; 
		rom[ 305  ] = 0; 
		rom[ 306  ] = 0; 
		rom[ 307  ] = 0; 
		rom[ 308  ] = 0; 
		rom[ 309  ] = 0; 
		rom[ 310  ] = 0; 
		rom[ 311  ] = 0; 
		rom[ 312  ] = 0; 
		rom[ 313  ] = 0; 
		rom[ 314  ] = 0; 
		rom[ 315  ] = 0; 
		rom[ 316  ] = 0; 
		rom[ 317  ] = 8192; 
		rom[ 318  ] = 8192; 
		rom[ 319  ] = 8192; 
		rom[ 320  ] = 0; 
		rom[ 321  ] = 0; 
		rom[ 322  ] = 0; 
		rom[ 323  ] = 0; 
		rom[ 324  ] = 0; 
		rom[ 325  ] = 0; 
		rom[ 326  ] = 0; 
		rom[ 327  ] = 8192; 
		rom[ 328  ] = 0; 
		rom[ 329  ] = 0; 
		rom[ 330  ] = 0; 
		rom[ 331  ] = 0; 
		rom[ 332  ] = 0; 
		rom[ 333  ] = 0; 
		rom[ 334  ] = 0; 
		rom[ 335  ] = 0; 
		rom[ 336  ] = 8192; 
		rom[ 337  ] = 8192; 
		rom[ 338  ] = 0; 
		rom[ 339  ] = 0; 
		rom[ 340  ] = 0; 
		rom[ 341  ] = 0; 
		rom[ 342  ] = 0; 
		rom[ 343  ] = 0; 
		rom[ 344  ] = 0; 
		rom[ 345  ] = 0; 
		rom[ 346  ] = 0; 
		rom[ 347  ] = 0; 
		rom[ 348  ] = 0; 
		rom[ 349  ] = 0; 
		rom[ 350  ] = 0; 
		rom[ 351  ] = 0; 
		rom[ 352  ] = 0; 
		rom[ 353  ] = 0; 
		rom[ 354  ] = 0; 
		rom[ 355  ] = 0; 
		rom[ 356  ] = 0; 
		rom[ 357  ] = 0; 
		rom[ 358  ] = 0; 
		rom[ 359  ] = 8192; 
		rom[ 360  ] = 8192; 
		rom[ 361  ] = 8192; 
		rom[ 362  ] = 8192; 
		rom[ 363  ] = 8192; 
		rom[ 364  ] = 0; 
		rom[ 365  ] = 0; 
		rom[ 366  ] = 8192; 
		rom[ 367  ] = 8192; 
		rom[ 368  ] = 0; 
		rom[ 369  ] = 0; 
		rom[ 370  ] = 0; 
		rom[ 371  ] = 0; 
		rom[ 372  ] = 0; 
		rom[ 373  ] = 8192; 
		rom[ 374  ] = 8192; 
		rom[ 375  ] = 8192; 
		rom[ 376  ] = 0; 
		rom[ 377  ] = 0; 
		rom[ 378  ] = 0; 
		rom[ 379  ] = 0; 
		rom[ 380  ] = 0; 
		rom[ 381  ] = 0; 
		rom[ 382  ] = 0; 
		rom[ 383  ] = 0; 
		rom[ 384  ] = 0; 
		rom[ 385  ] = 0; 
		rom[ 386  ] = 0; 
		rom[ 387  ] = 0; 
		rom[ 388  ] = 0; 
		rom[ 389  ] = 0; 
		rom[ 390  ] = 0; 
		rom[ 391  ] = 0; 
		rom[ 392  ] = 0; 
		rom[ 393  ] = 0; 
		rom[ 394  ] = 0; 
		rom[ 395  ] = 0; 
		rom[ 396  ] = 0; 
		rom[ 397  ] = 0; 
		rom[ 398  ] = 0; 
		rom[ 399  ] = 0; 
		rom[ 400  ] = 0; 
		rom[ 401  ] = 0; 
		rom[ 402  ] = 0; 
		rom[ 403  ] = 0; 
		rom[ 404  ] = 0; 
		rom[ 405  ] = 0; 
		rom[ 406  ] = 0; 
		rom[ 407  ] = 0; 
		rom[ 408  ] = 0; 
		rom[ 409  ] = 0; 
		rom[ 410  ] = 0; 
		rom[ 411  ] = 0; 
		rom[ 412  ] = 8192; 
		rom[ 413  ] = 0; 
		rom[ 414  ] = 0; 
		rom[ 415  ] = 8192; 
		rom[ 416  ] = 8192; 
		rom[ 417  ] = 0; 
		rom[ 418  ] = 0; 
		rom[ 419  ] = 0; 
		rom[ 420  ] = 0; 
		rom[ 421  ] = 0; 
		rom[ 422  ] = 0; 
		rom[ 423  ] = 0; 
		rom[ 424  ] = 0; 
		rom[ 425  ] = 0; 
		rom[ 426  ] = 0; 
		rom[ 427  ] = 0; 
		rom[ 428  ] = 0; 
		rom[ 429  ] = 0; 
		rom[ 430  ] = 0; 
		rom[ 431  ] = 0; 
		rom[ 432  ] = 0; 
		rom[ 433  ] = 0; 
		rom[ 434  ] = 0; 
		rom[ 435  ] = 0; 
		rom[ 436  ] = 0; 
		rom[ 437  ] = 0; 
		rom[ 438  ] = 0; 
		rom[ 439  ] = 0; 
		rom[ 440  ] = 0; 
		rom[ 441  ] = 0; 
		rom[ 442  ] = 0; 
		rom[ 443  ] = 0; 
		rom[ 444  ] = 8192; 
		rom[ 445  ] = 0; 
		rom[ 446  ] = 0; 
		rom[ 447  ] = 0; 
		rom[ 448  ] = 0; 
		rom[ 449  ] = 0; 
		rom[ 450  ] = 0; 
		rom[ 451  ] = 8192; 
		rom[ 452  ] = 0; 
		rom[ 453  ] = 8192; 
		rom[ 454  ] = 8192; 
		rom[ 455  ] = 0; 
		rom[ 456  ] = 0; 
		rom[ 457  ] = 0; 
		rom[ 458  ] = 0; 
		rom[ 459  ] = 8192; 
		rom[ 460  ] = 8192; 
		rom[ 461  ] = 8192; 
		rom[ 462  ] = 0; 
		rom[ 463  ] = 8192; 
		rom[ 464  ] = 8192; 
		rom[ 465  ] = 0; 
		rom[ 466  ] = 0; 
		rom[ 467  ] = 0; 
		rom[ 468  ] = 0; 
		rom[ 469  ] = 0; 
		rom[ 470  ] = 0; 
		rom[ 471  ] = 0; 
		rom[ 472  ] = 0; 
		rom[ 473  ] = 8192; 
		rom[ 474  ] = 0; 
		rom[ 475  ] = 0; 
		rom[ 476  ] = 0; 
		rom[ 477  ] = 0; 
		rom[ 478  ] = 8192; 
		rom[ 479  ] = 0; 
		rom[ 480  ] = 0; 
		rom[ 481  ] = 8192; 
		rom[ 482  ] = 0; 
		rom[ 483  ] = 0; 
		rom[ 484  ] = 0; 
		rom[ 485  ] = 0; 
		rom[ 486  ] = 0; 
		rom[ 487  ] = 0; 
		rom[ 488  ] = 0; 
		rom[ 489  ] = 0; 
		rom[ 490  ] = 8192; 
		rom[ 491  ] = 0; 
		rom[ 492  ] = 0; 
		rom[ 493  ] = 0; 
		rom[ 494  ] = 0; 
		rom[ 495  ] = 0; 
		rom[ 496  ] = 0; 
		rom[ 497  ] = 0; 
		rom[ 498  ] = 0; 
		rom[ 499  ] = 0; 
		rom[ 500  ] = 0; 
		rom[ 501  ] = 0; 
		rom[ 502  ] = 0; 
		rom[ 503  ] = 0; 
		rom[ 504  ] = 0; 
		rom[ 505  ] = 0; 
		rom[ 506  ] = 0; 
		rom[ 507  ] = 0; 
		rom[ 508  ] = 0; 
		rom[ 509  ] = 0; 
		rom[ 510  ] = 0; 
		rom[ 511  ] = 0; 
		rom[ 512  ] = 0; 
		rom[ 513  ] = 0; 
		rom[ 514  ] = 0; 
		rom[ 515  ] = 0; 
		rom[ 516  ] = 0; 
		rom[ 517  ] = 0; 
		rom[ 518  ] = 0; 
		rom[ 519  ] = 0; 
		rom[ 520  ] = 8192; 
		rom[ 521  ] = 8192; 
		rom[ 522  ] = 0; 
		rom[ 523  ] = 0; 
		rom[ 524  ] = 0; 
		rom[ 525  ] = 8192; 
		rom[ 526  ] = 0; 
		rom[ 527  ] = 0; 
		rom[ 528  ] = 0; 
		rom[ 529  ] = 8192; 
		rom[ 530  ] = 0; 
		rom[ 531  ] = 0; 
		rom[ 532  ] = 0; 
		rom[ 533  ] = 0; 
		rom[ 534  ] = 0; 
		rom[ 535  ] = 0; 
		rom[ 536  ] = 0; 
		rom[ 537  ] = 0; 
		rom[ 538  ] = 0; 
		rom[ 539  ] = 0; 
		rom[ 540  ] = 0; 
		rom[ 541  ] = 0; 
		rom[ 542  ] = 8192; 
		rom[ 543  ] = 0; 
		rom[ 544  ] = 0; 
		rom[ 545  ] = 0; 
		rom[ 546  ] = 8192; 
		rom[ 547  ] = 0; 
		rom[ 548  ] = 8192; 
		rom[ 549  ] = 8192; 
		rom[ 550  ] = 0; 
		rom[ 551  ] = 0; 
		rom[ 552  ] = 0; 
		rom[ 553  ] = 0; 
		rom[ 554  ] = 8192; 
		rom[ 555  ] = 0; 
		rom[ 556  ] = 0; 
		rom[ 557  ] = 0; 
		rom[ 558  ] = 0; 
		rom[ 559  ] = 8192; 
		rom[ 560  ] = 0; 
		rom[ 561  ] = 0; 
		rom[ 562  ] = 0; 
		rom[ 563  ] = 0; 
		rom[ 564  ] = 0; 
		rom[ 565  ] = 0; 
		rom[ 566  ] = 0; 
		rom[ 567  ] = 0; 
		rom[ 568  ] = 0; 
		rom[ 569  ] = 0; 
		rom[ 570  ] = 0; 
		rom[ 571  ] = 0; 
		rom[ 572  ] = 0; 
		rom[ 573  ] = 0; 
		rom[ 574  ] = 0; 
		rom[ 575  ] = 0; 
		rom[ 576  ] = 0; 
		rom[ 577  ] = 0; 
		rom[ 578  ] = 0; 
		rom[ 579  ] = 0; 
		rom[ 580  ] = 0; 
		rom[ 581  ] = 0; 
		rom[ 582  ] = 0; 
		rom[ 583  ] = 0; 
		rom[ 584  ] = 0; 
		rom[ 585  ] = 0; 
		rom[ 586  ] = 0; 
		rom[ 587  ] = 8192; 
		rom[ 588  ] = 8192; 
		rom[ 589  ] = 0; 
		rom[ 590  ] = 0; 
		rom[ 591  ] = 8192; 
		rom[ 592  ] = 8192; 
		rom[ 593  ] = 0; 
		rom[ 594  ] = 8192; 
		rom[ 595  ] = 8192; 
		rom[ 596  ] = 0; 
		rom[ 597  ] = 0; 
		rom[ 598  ] = 0; 
		rom[ 599  ] = 0; 
		rom[ 600  ] = 0; 
		rom[ 601  ] = 0; 
		rom[ 602  ] = 0; 
		rom[ 603  ] = 0; 
		rom[ 604  ] = 0; 
		rom[ 605  ] = 0; 
		rom[ 606  ] = 0; 
		rom[ 607  ] = 0; 
		rom[ 608  ] = 0; 
		rom[ 609  ] = 0; 
		rom[ 610  ] = 0; 
		rom[ 611  ] = 0; 
		rom[ 612  ] = 0; 
		rom[ 613  ] = 0; 
		rom[ 614  ] = 0; 
		rom[ 615  ] = 0; 
		rom[ 616  ] = 0; 
		rom[ 617  ] = 0; 
		rom[ 618  ] = 0; 
		rom[ 619  ] = 0; 
		rom[ 620  ] = 0; 
		rom[ 621  ] = 0; 
		rom[ 622  ] = 0; 
		rom[ 623  ] = 0; 
		rom[ 624  ] = 8192; 
		rom[ 625  ] = 8192; 
		rom[ 626  ] = 0; 
		rom[ 627  ] = 0; 
		rom[ 628  ] = 0; 
		rom[ 629  ] = 0; 
		rom[ 630  ] = 0; 
		rom[ 631  ] = 0; 
		rom[ 632  ] = 0; 
		rom[ 633  ] = 0; 
		rom[ 634  ] = 0; 
		rom[ 635  ] = 0; 
		rom[ 636  ] = 0; 
		rom[ 637  ] = 0; 
		rom[ 638  ] = 0; 
		rom[ 639  ] = 0; 
		rom[ 640  ] = 0; 
		rom[ 641  ] = 0; 
		rom[ 642  ] = 0; 
		rom[ 643  ] = 0; 
		rom[ 644  ] = 0; 
		rom[ 645  ] = 0; 
		rom[ 646  ] = 0; 
		rom[ 647  ] = 0; 
		rom[ 648  ] = 0; 
		rom[ 649  ] = 0; 
		rom[ 650  ] = 0; 
		rom[ 651  ] = 0; 
		rom[ 652  ] = 0; 
		rom[ 653  ] = 0; 
		rom[ 654  ] = 0; 
		rom[ 655  ] = 8192; 
		rom[ 656  ] = 0; 
		rom[ 657  ] = 0; 
		rom[ 658  ] = 0; 
		rom[ 659  ] = 8192; 
		rom[ 660  ] = 0; 
		rom[ 661  ] = 0; 
		rom[ 662  ] = 0; 
		rom[ 663  ] = 0; 
		rom[ 664  ] = 0; 
		rom[ 665  ] = 8192; 
		rom[ 666  ] = 8192; 
		rom[ 667  ] = 0; 
		rom[ 668  ] = 0; 
		rom[ 669  ] = 0; 
		rom[ 670  ] = 0; 
		rom[ 671  ] = 0; 
		rom[ 672  ] = 0; 
		rom[ 673  ] = 0; 
		rom[ 674  ] = 0; 
		rom[ 675  ] = 8192; 
		rom[ 676  ] = 0; 
		rom[ 677  ] = 0; 
		rom[ 678  ] = 8192; 
		rom[ 679  ] = 8192; 
		rom[ 680  ] = 8192; 
		rom[ 681  ] = 0; 
		rom[ 682  ] = 0; 
		rom[ 683  ] = 8192; 
		rom[ 684  ] = 0; 
		rom[ 685  ] = 0; 
		rom[ 686  ] = 8192; 
		rom[ 687  ] = 0; 
		rom[ 688  ] = 0; 
		rom[ 689  ] = 0; 
		rom[ 690  ] = 0; 
		rom[ 691  ] = 8192; 
		rom[ 692  ] = 0; 
		rom[ 693  ] = 0; 
		rom[ 694  ] = 8192; 
		rom[ 695  ] = 0; 
		rom[ 696  ] = 0; 
		rom[ 697  ] = 0; 
		rom[ 698  ] = 0; 
		rom[ 699  ] = 8192; 
		rom[ 700  ] = 8192; 
		rom[ 701  ] = 0; 
		rom[ 702  ] = 0; 
		rom[ 703  ] = 0; 
		rom[ 704  ] = 8192; 
		rom[ 705  ] = 8192; 
		rom[ 706  ] = 8192; 
		rom[ 707  ] = 0; 
		rom[ 708  ] = 0; 
		rom[ 709  ] = 0; 
		rom[ 710  ] = 0; 
		rom[ 711  ] = 0; 
		rom[ 712  ] = 0; 
		rom[ 713  ] = 0; 
		rom[ 714  ] = 0; 
		rom[ 715  ] = 0; 
		rom[ 716  ] = 0; 
		rom[ 717  ] = 0; 
		rom[ 718  ] = 0; 
		rom[ 719  ] = 0; 
		rom[ 720  ] = 0; 
		rom[ 721  ] = 0; 
		rom[ 722  ] = 8192; 
		rom[ 723  ] = 0; 
		rom[ 724  ] = 0; 
		rom[ 725  ] = 0; 
		rom[ 726  ] = 8192; 
		rom[ 727  ] = 0; 
		rom[ 728  ] = 0; 
		rom[ 729  ] = 0; 
		rom[ 730  ] = 0; 
		rom[ 731  ] = 0; 
		rom[ 732  ] = 0; 
		rom[ 733  ] = 0; 
		rom[ 734  ] = 0; 
		rom[ 735  ] = 0; 
		rom[ 736  ] = 0; 
		rom[ 737  ] = 0; 
		rom[ 738  ] = 0; 
		rom[ 739  ] = 0; 
		rom[ 740  ] = 0; 
		rom[ 741  ] = 0; 
		rom[ 742  ] = 0; 
		rom[ 743  ] = 0; 
		rom[ 744  ] = 0; 
		rom[ 745  ] = 0; 
		rom[ 746  ] = 0; 
		rom[ 747  ] = 0; 
		rom[ 748  ] = 0; 
		rom[ 749  ] = 0; 
		rom[ 750  ] = 0; 
		rom[ 751  ] = 8192; 
		rom[ 752  ] = 8192; 
		rom[ 753  ] = 0; 
		rom[ 754  ] = 0; 
		rom[ 755  ] = 0; 
		rom[ 756  ] = 8192; 
		rom[ 757  ] = 8192; 
		rom[ 758  ] = 8192; 
		rom[ 759  ] = 0; 
		rom[ 760  ] = 0; 
		rom[ 761  ] = 8192; 
		rom[ 762  ] = 0; 
		rom[ 763  ] = 0; 
		rom[ 764  ] = 0; 
		rom[ 765  ] = 0; 
		rom[ 766  ] = 0; 
		rom[ 767  ] = 0; 
		rom[ 768  ] = 0; 
		rom[ 769  ] = 0; 
		rom[ 770  ] = 8192; 
		rom[ 771  ] = 0; 
		rom[ 772  ] = 0; 
		rom[ 773  ] = 0; 
		rom[ 774  ] = 0; 
		rom[ 775  ] = 8192; 
		rom[ 776  ] = 0; 
		rom[ 777  ] = 0; 
		rom[ 778  ] = 8192; 
		rom[ 779  ] = 0; 
		rom[ 780  ] = 0; 
		rom[ 781  ] = 0; 
		rom[ 782  ] = 0; 
		rom[ 783  ] = 0; 
		rom[ 784  ] = 8192; 
		rom[ 785  ] = 0; 
		rom[ 786  ] = 8192; 
		rom[ 787  ] = 0; 
		rom[ 788  ] = 0; 
		rom[ 789  ] = 0; 
		rom[ 790  ] = 0; 
		rom[ 791  ] = 0; 
		rom[ 792  ] = 0; 
		rom[ 793  ] = 0; 
		rom[ 794  ] = 0; 
		rom[ 795  ] = 0; 
		rom[ 796  ] = 0; 
		rom[ 797  ] = 0; 
		rom[ 798  ] = 0; 
		rom[ 799  ] = 0; 
		rom[ 800  ] = 8192; 
		rom[ 801  ] = 0; 
		rom[ 802  ] = 0; 
		rom[ 803  ] = 0; 
		rom[ 804  ] = 0; 
		rom[ 805  ] = 0; 
		rom[ 806  ] = 0; 
		rom[ 807  ] = 8192; 
		rom[ 808  ] = 0; 
		rom[ 809  ] = 0; 
		rom[ 810  ] = 0; 
		rom[ 811  ] = 0; 
		rom[ 812  ] = 0; 
		rom[ 813  ] = 0; 
		rom[ 814  ] = 0; 
		rom[ 815  ] = 0; 
		rom[ 816  ] = 0; 
		rom[ 817  ] = 0; 
		rom[ 818  ] = 0; 
		rom[ 819  ] = 8192; 
		rom[ 820  ] = 0; 
		rom[ 821  ] = 0; 
		rom[ 822  ] = 0; 
		rom[ 823  ] = 0; 
		rom[ 824  ] = 0; 
		rom[ 825  ] = 0; 
		rom[ 826  ] = 0; 
		rom[ 827  ] = 0; 
		rom[ 828  ] = 0; 
		rom[ 829  ] = 0; 
		rom[ 830  ] = 0; 
		rom[ 831  ] = 0; 
		rom[ 832  ] = 0; 
		rom[ 833  ] = 8192; 
		rom[ 834  ] = 0; 
		rom[ 835  ] = 0; 
		rom[ 836  ] = 0; 
		rom[ 837  ] = 0; 
		rom[ 838  ] = 0; 
		rom[ 839  ] = 0; 
		rom[ 840  ] = 0; 
		rom[ 841  ] = 0; 
		rom[ 842  ] = 0; 
		rom[ 843  ] = 0; 
		rom[ 844  ] = 0; 
		rom[ 845  ] = 0; 
		rom[ 846  ] = 0; 
		rom[ 847  ] = 0; 
		rom[ 848  ] = 0; 
		rom[ 849  ] = 0; 
		rom[ 850  ] = 0; 
		rom[ 851  ] = 8192; 
		rom[ 852  ] = 0; 
		rom[ 853  ] = 0; 
		rom[ 854  ] = 0; 
		rom[ 855  ] = 8192; 
		rom[ 856  ] = 0; 
		rom[ 857  ] = 0; 
		rom[ 858  ] = 0; 
		rom[ 859  ] = 8192; 
		rom[ 860  ] = 0; 
		rom[ 861  ] = 8192; 
		rom[ 862  ] = 8192; 
		rom[ 863  ] = 0; 
		rom[ 864  ] = 0; 
		rom[ 865  ] = 8192; 
		rom[ 866  ] = 8192; 
		rom[ 867  ] = 0; 
		rom[ 868  ] = 8192; 
		rom[ 869  ] = 0; 
		rom[ 870  ] = 0; 
		rom[ 871  ] = 0; 
		rom[ 872  ] = 0; 
		rom[ 873  ] = 0; 
		rom[ 874  ] = 0; 
		rom[ 875  ] = 0; 
		rom[ 876  ] = 8192; 
		rom[ 877  ] = 0; 
		rom[ 878  ] = 0; 
		rom[ 879  ] = 0; 
		rom[ 880  ] = 0; 
		rom[ 881  ] = 0; 
		rom[ 882  ] = 0; 
		rom[ 883  ] = 0; 
		rom[ 884  ] = 0; 
		rom[ 885  ] = 0; 
		rom[ 886  ] = 0; 
		rom[ 887  ] = 0; 
		rom[ 888  ] = 0; 
		rom[ 889  ] = 0; 
		rom[ 890  ] = 0; 
		rom[ 891  ] = 0; 
		rom[ 892  ] = 0; 
		rom[ 893  ] = 0; 
		rom[ 894  ] = 0; 
		rom[ 895  ] = 0; 
		rom[ 896  ] = 0; 
		rom[ 897  ] = 0; 
		rom[ 898  ] = 0; 
		rom[ 899  ] = 0; 
		rom[ 900  ] = 0; 
		rom[ 901  ] = 0; 
		rom[ 902  ] = 0; 
		rom[ 903  ] = 0; 
		rom[ 904  ] = 0; 
		rom[ 905  ] = 0; 
		rom[ 906  ] = 0; 
		rom[ 907  ] = 0; 
		rom[ 908  ] = 0; 
		rom[ 909  ] = 0; 
		rom[ 910  ] = 0; 
		rom[ 911  ] = 8192; 
		rom[ 912  ] = 8192; 
		rom[ 913  ] = 0; 
		rom[ 914  ] = 0; 
		rom[ 915  ] = 0; 
		rom[ 916  ] = 0; 
		rom[ 917  ] = 0; 
		rom[ 918  ] = 0; 
		rom[ 919  ] = 0; 
		rom[ 920  ] = 8192; 
		rom[ 921  ] = 0; 
		rom[ 922  ] = 0; 
		rom[ 923  ] = 0; 
		rom[ 924  ] = 0; 
		rom[ 925  ] = 0; 
		rom[ 926  ] = 0; 
		rom[ 927  ] = 0; 
		rom[ 928  ] = 0; 
		rom[ 929  ] = 0; 
		rom[ 930  ] = 0; 
		rom[ 931  ] = 0; 
		rom[ 932  ] = 0; 
		rom[ 933  ] = 0; 
		rom[ 934  ] = 0; 
		rom[ 935  ] = 0; 
		rom[ 936  ] = 0; 
		rom[ 937  ] = 0; 
		rom[ 938  ] = 0; 
		rom[ 939  ] = 0; 
		rom[ 940  ] = 0; 
		rom[ 941  ] = 0; 
		rom[ 942  ] = 0; 
		rom[ 943  ] = 0; 
		rom[ 944  ] = 0; 
		rom[ 945  ] = 0; 
		rom[ 946  ] = 8192; 
		rom[ 947  ] = 8192; 
		rom[ 948  ] = 0; 
		rom[ 949  ] = 8192; 
		rom[ 950  ] = 8192; 
		rom[ 951  ] = 8192; 
		rom[ 952  ] = 0; 
		rom[ 953  ] = 8192; 
		rom[ 954  ] = 0; 
		rom[ 955  ] = 8192; 
		rom[ 956  ] = 0; 
		rom[ 957  ] = 8192; 
		rom[ 958  ] = 0; 
		rom[ 959  ] = 8192; 
		rom[ 960  ] = 0; 
		rom[ 961  ] = 0; 
		rom[ 962  ] = 8192; 
		rom[ 963  ] = 0; 
		rom[ 964  ] = 0; 
		rom[ 965  ] = 8192; 
		rom[ 966  ] = 8192; 
		rom[ 967  ] = 0; 
		rom[ 968  ] = 8192; 
		rom[ 969  ] = 0; 
		rom[ 970  ] = 0; 
		rom[ 971  ] = 0; 
		rom[ 972  ] = 0; 
		rom[ 973  ] = 0; 
		rom[ 974  ] = 0; 
		rom[ 975  ] = 0; 
		rom[ 976  ] = 0; 
		rom[ 977  ] = 8192; 
		rom[ 978  ] = 8192; 
		rom[ 979  ] = 0; 
		rom[ 980  ] = 8192; 
		rom[ 981  ] = 8192; 
		rom[ 982  ] = 0; 
		rom[ 983  ] = 0; 
		rom[ 984  ] = 0; 
		rom[ 985  ] = 0; 
		rom[ 986  ] = 0; 
		rom[ 987  ] = 0; 
		rom[ 988  ] = 0; 
		rom[ 989  ] = 0; 
		rom[ 990  ] = 8192; 
		rom[ 991  ] = 8192; 
		rom[ 992  ] = 0; 
		rom[ 993  ] = 0; 
		rom[ 994  ] = 0; 
		rom[ 995  ] = 0; 
		rom[ 996  ] = 0; 
		rom[ 997  ] = 0; 
		rom[ 998  ] = 0; 
		rom[ 999  ] = 0; 
		rom[ 1000 ] = 0; 
		rom[ 1001 ] = 0; 
		rom[ 1002 ] = 0; 
		rom[ 1003 ] = 0; 
		rom[ 1004 ] = 0; 
		rom[ 1005 ] = 0; 
		rom[ 1006 ] = 0; 
		rom[ 1007 ] = 0; 
		rom[ 1008 ] = 0; 
		rom[ 1009 ] = 8192; 
		rom[ 1010 ] = 0; 
		rom[ 1011 ] = 0; 
		rom[ 1012 ] = 8192; 
		rom[ 1013 ] = 8192; 
		rom[ 1014 ] = 0; 
		rom[ 1015 ] = 0; 
		rom[ 1016 ] = 8192; 
		rom[ 1017 ] = 8192; 
		rom[ 1018 ] = 8192; 
		rom[ 1019 ] = 0; 
		rom[ 1020 ] = 0; 
		rom[ 1021 ] = 8192; 
		rom[ 1022 ] = 0; 
		rom[ 1023 ] = 0; 
		rom[ 1024 ] = 0; 
		rom[ 1025 ] = 0; 
		rom[ 1026 ] = 0; 
		rom[ 1027 ] = 0; 
		rom[ 1028 ] = 0; 
		rom[ 1029 ] = 0; 
		rom[ 1030 ] = 0; 
		rom[ 1031 ] = 0; 
		rom[ 1032 ] = 0; 
		rom[ 1033 ] = 0; 
		rom[ 1034 ] = 0; 
		rom[ 1035 ] = 0; 
		rom[ 1036 ] = 0; 
		rom[ 1037 ] = 0; 
		rom[ 1038 ] = 0; 
		rom[ 1039 ] = 0; 
		rom[ 1040 ] = 0; 
		rom[ 1041 ] = 0; 
		rom[ 1042 ] = 0; 
		rom[ 1043 ] = 0; 
		rom[ 1044 ] = 8192; 
		rom[ 1045 ] = 0; 
		rom[ 1046 ] = 8192; 
		rom[ 1047 ] = 8192; 
		rom[ 1048 ] = 0; 
		rom[ 1049 ] = 0; 
		rom[ 1050 ] = 0; 
		rom[ 1051 ] = 0; 
		rom[ 1052 ] = 0; 
		rom[ 1053 ] = 0; 
		rom[ 1054 ] = 0; 
		rom[ 1055 ] = 0; 
		rom[ 1056 ] = 0; 
		rom[ 1057 ] = 8192; 
		rom[ 1058 ] = 8192; 
		rom[ 1059 ] = 0; 
		rom[ 1060 ] = 0; 
		rom[ 1061 ] = 0; 
		rom[ 1062 ] = 0; 
		rom[ 1063 ] = 0; 
		rom[ 1064 ] = 0; 
		rom[ 1065 ] = 0; 
		rom[ 1066 ] = 0; 
		rom[ 1067 ] = 0; 
		rom[ 1068 ] = 0; 
		rom[ 1069 ] = 0; 
		rom[ 1070 ] = 0; 
		rom[ 1071 ] = 0; 
		rom[ 1072 ] = 0; 
		rom[ 1073 ] = 0; 
		rom[ 1074 ] = 8192; 
		rom[ 1075 ] = 0; 
		rom[ 1076 ] = 0; 
		rom[ 1077 ] = 0; 
		rom[ 1078 ] = 0; 
		rom[ 1079 ] = 0; 
		rom[ 1080 ] = 8192; 
		rom[ 1081 ] = 8192; 
		rom[ 1082 ] = 0; 
		rom[ 1083 ] = 8192; 
		rom[ 1084 ] = 0; 
		rom[ 1085 ] = 0; 
		rom[ 1086 ] = 0; 
		rom[ 1087 ] = 8192; 
		rom[ 1088 ] = 0; 
		rom[ 1089 ] = 0; 
		rom[ 1090 ] = 0; 
		rom[ 1091 ] = 0; 
		rom[ 1092 ] = 0; 
		rom[ 1093 ] = 0; 
		rom[ 1094 ] = 8192; 
		rom[ 1095 ] = 8192; 
		rom[ 1096 ] = 8192; 
		rom[ 1097 ] = 0; 
		rom[ 1098 ] = 8192; 
		rom[ 1099 ] = 0; 
		rom[ 1100 ] = 8192; 
		rom[ 1101 ] = 0; 
		rom[ 1102 ] = 0; 
		rom[ 1103 ] = 0; 
		rom[ 1104 ] = 0; 
		rom[ 1105 ] = 0; 
		rom[ 1106 ] = 0; 
		rom[ 1107 ] = 0; 
		rom[ 1108 ] = 0; 
		rom[ 1109 ] = 0; 
		rom[ 1110 ] = 0; 
		rom[ 1111 ] = 0; 
		rom[ 1112 ] = 0; 
		rom[ 1113 ] = 0; 
		rom[ 1114 ] = 0; 
		rom[ 1115 ] = 0; 
		rom[ 1116 ] = 0; 
		rom[ 1117 ] = 0; 
		rom[ 1118 ] = 0; 
		rom[ 1119 ] = 0; 
		rom[ 1120 ] = 0; 
		rom[ 1121 ] = 0; 
		rom[ 1122 ] = 0; 
		rom[ 1123 ] = 0; 
		rom[ 1124 ] = 0; 
		rom[ 1125 ] = 0; 
		rom[ 1126 ] = 0; 
		rom[ 1127 ] = 0; 
		rom[ 1128 ] = 0; 
		rom[ 1129 ] = 0; 
		rom[ 1130 ] = 0; 
		rom[ 1131 ] = 0; 
		rom[ 1132 ] = 0; 
		rom[ 1133 ] = 0; 
		rom[ 1134 ] = 0; 
		rom[ 1135 ] = 0; 
		rom[ 1136 ] = 0; 
		rom[ 1137 ] = 8192; 
		rom[ 1138 ] = 8192; 
		rom[ 1139 ] = 8192; 
		rom[ 1140 ] = 0; 
		rom[ 1141 ] = 8192; 
		rom[ 1142 ] = 0; 
		rom[ 1143 ] = 0; 
		rom[ 1144 ] = 0; 
		rom[ 1145 ] = 0; 
		rom[ 1146 ] = 0; 
		rom[ 1147 ] = 0; 
		rom[ 1148 ] = 0; 
		rom[ 1149 ] = 0; 
		rom[ 1150 ] = 0; 
		rom[ 1151 ] = 0; 
		rom[ 1152 ] = 0; 
		rom[ 1153 ] = 0; 
		rom[ 1154 ] = 0; 
		rom[ 1155 ] = 0; 
		rom[ 1156 ] = 0; 
		rom[ 1157 ] = 0; 
		rom[ 1158 ] = 0; 
		rom[ 1159 ] = 0; 
		rom[ 1160 ] = 0; 
		rom[ 1161 ] = 8192; 
		rom[ 1162 ] = 0; 
		rom[ 1163 ] = 0; 
		rom[ 1164 ] = 0; 
		rom[ 1165 ] = 0; 
		rom[ 1166 ] = 0; 
		rom[ 1167 ] = 0; 
		rom[ 1168 ] = 0; 
		rom[ 1169 ] = 0; 
		rom[ 1170 ] = 0; 
		rom[ 1171 ] = 0; 
		rom[ 1172 ] = 0; 
		rom[ 1173 ] = 0; 
		rom[ 1174 ] = 0; 
		rom[ 1175 ] = 0; 
		rom[ 1176 ] = 0; 
		rom[ 1177 ] = 8192; 
		rom[ 1178 ] = 0; 
		rom[ 1179 ] = 8192; 
		rom[ 1180 ] = 8192; 
		rom[ 1181 ] = 8192; 
		rom[ 1182 ] = 0; 
		rom[ 1183 ] = 0; 
		rom[ 1184 ] = 8192; 
		rom[ 1185 ] = 0; 
		rom[ 1186 ] = 0; 
		rom[ 1187 ] = 0; 
		rom[ 1188 ] = 0; 
		rom[ 1189 ] = 0; 
		rom[ 1190 ] = 0; 
		rom[ 1191 ] = 0; 
		rom[ 1192 ] = 0; 
		rom[ 1193 ] = 0; 
		rom[ 1194 ] = 0; 
		rom[ 1195 ] = 0; 
		rom[ 1196 ] = 0; 
		rom[ 1197 ] = 0; 
		rom[ 1198 ] = 0; 
		rom[ 1199 ] = 0; 
		rom[ 1200 ] = 0; 
		rom[ 1201 ] = 0; 
		rom[ 1202 ] = 0; 
		rom[ 1203 ] = 0; 
		rom[ 1204 ] = 0; 
		rom[ 1205 ] = 0; 
		rom[ 1206 ] = 0; 
		rom[ 1207 ] = 0; 
		rom[ 1208 ] = 0; 
		rom[ 1209 ] = 8192; 
		rom[ 1210 ] = 8192; 
		rom[ 1211 ] = 8192; 
		rom[ 1212 ] = 8192; 
		rom[ 1213 ] = 0; 
		rom[ 1214 ] = 0; 
		rom[ 1215 ] = 0; 
		rom[ 1216 ] = 0; 
		rom[ 1217 ] = 0; 
		rom[ 1218 ] = 0; 
		rom[ 1219 ] = 0; 
		rom[ 1220 ] = 0; 
		rom[ 1221 ] = 0; 
		rom[ 1222 ] = 0; 
		rom[ 1223 ] = 0; 
		rom[ 1224 ] = 0; 
		rom[ 1225 ] = 0; 
		rom[ 1226 ] = 8192; 
		rom[ 1227 ] = 0; 
		rom[ 1228 ] = 0; 
		rom[ 1229 ] = 0; 
		rom[ 1230 ] = 0; 
		rom[ 1231 ] = 0; 
		rom[ 1232 ] = 0; 
		rom[ 1233 ] = 8192; 
		rom[ 1234 ] = 8192; 
		rom[ 1235 ] = 0; 
		rom[ 1236 ] = 0; 
		rom[ 1237 ] = 0; 
		rom[ 1238 ] = 8192; 
		rom[ 1239 ] = 0; 
		rom[ 1240 ] = 0; 
		rom[ 1241 ] = 0; 
		rom[ 1242 ] = 0; 
		rom[ 1243 ] = 8192; 
		rom[ 1244 ] = 0; 
		rom[ 1245 ] = 0; 
		rom[ 1246 ] = 0; 
		rom[ 1247 ] = 0; 
		rom[ 1248 ] = 0; 
		rom[ 1249 ] = 0; 
		rom[ 1250 ] = 0; 
		rom[ 1251 ] = 0; 
		rom[ 1252 ] = 0; 
		rom[ 1253 ] = 0; 
		rom[ 1254 ] = 0; 
		rom[ 1255 ] = 0; 
		rom[ 1256 ] = 8192; 
		rom[ 1257 ] = 0; 
		rom[ 1258 ] = 0; 
		rom[ 1259 ] = 0; 
		rom[ 1260 ] = 0; 
		rom[ 1261 ] = 0; 
		rom[ 1262 ] = 8192; 
		rom[ 1263 ] = 0; 
		rom[ 1264 ] = 8192; 
		rom[ 1265 ] = 8192; 
		rom[ 1266 ] = 8192; 
		rom[ 1267 ] = 0; 
		rom[ 1268 ] = 0; 
		rom[ 1269 ] = 0; 
		rom[ 1270 ] = 0; 
		rom[ 1271 ] = 0; 
		rom[ 1272 ] = 0; 
		rom[ 1273 ] = 0; 
		rom[ 1274 ] = 0; 
		rom[ 1275 ] = 0; 
		rom[ 1276 ] = 0; 
		rom[ 1277 ] = 0; 
		rom[ 1278 ] = 0; 
		rom[ 1279 ] = 0; 
		rom[ 1280 ] = 0; 
		rom[ 1281 ] = 0; 
		rom[ 1282 ] = 0; 
		rom[ 1283 ] = 0; 
		rom[ 1284 ] = 0; 
		rom[ 1285 ] = 0; 
		rom[ 1286 ] = 0; 
		rom[ 1287 ] = 0; 
		rom[ 1288 ] = 0; 
		rom[ 1289 ] = 8192; 
		rom[ 1290 ] = 0; 
		rom[ 1291 ] = 8192; 
		rom[ 1292 ] = 0; 
		rom[ 1293 ] = 8192; 
		rom[ 1294 ] = 0; 
		rom[ 1295 ] = 8192; 
		rom[ 1296 ] = 0; 
		rom[ 1297 ] = 8192; 
		rom[ 1298 ] = 8192; 
		rom[ 1299 ] = 8192; 
		rom[ 1300 ] = 0; 
		rom[ 1301 ] = 8192; 
		rom[ 1302 ] = 8192; 
		rom[ 1303 ] = 8192; 
		rom[ 1304 ] = 8192; 
		rom[ 1305 ] = 8192; 
		rom[ 1306 ] = 8192; 
		rom[ 1307 ] = 8192; 
		rom[ 1308 ] = 8192; 
		rom[ 1309 ] = 0; 
		rom[ 1310 ] = 0; 
		rom[ 1311 ] = 0; 
		rom[ 1312 ] = 8192; 
		rom[ 1313 ] = 0; 
		rom[ 1314 ] = 0; 
		rom[ 1315 ] = 8192; 
		rom[ 1316 ] = 0; 
		rom[ 1317 ] = 0; 
		rom[ 1318 ] = 0; 
		rom[ 1319 ] = 0; 
		rom[ 1320 ] = 0; 
		rom[ 1321 ] = 0; 
		rom[ 1322 ] = 0; 
		rom[ 1323 ] = 0; 
		rom[ 1324 ] = 0; 
		rom[ 1325 ] = 8192; 
		rom[ 1326 ] = 8192; 
		rom[ 1327 ] = 0; 
		rom[ 1328 ] = 0; 
		rom[ 1329 ] = 8192; 
		rom[ 1330 ] = 8192; 
		rom[ 1331 ] = 0; 
		rom[ 1332 ] = 0; 
		rom[ 1333 ] = 0; 
		rom[ 1334 ] = 0; 
		rom[ 1335 ] = 8192; 
		rom[ 1336 ] = 8192; 
		rom[ 1337 ] = 0; 
		rom[ 1338 ] = 0; 
		rom[ 1339 ] = 0; 
		rom[ 1340 ] = 0; 
		rom[ 1341 ] = 0; 
		rom[ 1342 ] = 0; 
		rom[ 1343 ] = 0; 
		rom[ 1344 ] = 0; 
		rom[ 1345 ] = 0; 
		rom[ 1346 ] = 0; 
		rom[ 1347 ] = 0; 
		rom[ 1348 ] = 8192; 
		rom[ 1349 ] = 0; 
		rom[ 1350 ] = 0; 
		rom[ 1351 ] = 0; 
		rom[ 1352 ] = 0; 
		rom[ 1353 ] = 8192; 
		rom[ 1354 ] = 8192; 
		rom[ 1355 ] = 8192; 
		rom[ 1356 ] = 0; 
		rom[ 1357 ] = 0; 
		rom[ 1358 ] = 0; 
		rom[ 1359 ] = 0; 
		rom[ 1360 ] = 0; 
		rom[ 1361 ] = 0; 
		rom[ 1362 ] = 0; 
		rom[ 1363 ] = 0; 
		rom[ 1364 ] = 0; 
		rom[ 1365 ] = 0; 
		rom[ 1366 ] = 0; 
		rom[ 1367 ] = 0; 
		rom[ 1368 ] = 0; 
		rom[ 1369 ] = 0; 
		rom[ 1370 ] = 8192; 
		rom[ 1371 ] = 8192; 
		rom[ 1372 ] = 8192; 
		rom[ 1373 ] = 0; 
		rom[ 1374 ] = 0; 
		rom[ 1375 ] = 0; 
		rom[ 1376 ] = 0; 
		rom[ 1377 ] = 8192; 
		rom[ 1378 ] = 0; 
		rom[ 1379 ] = 0; 
		rom[ 1380 ] = 0; 
		rom[ 1381 ] = 0; 
		rom[ 1382 ] = 0; 
		rom[ 1383 ] = 0; 
		rom[ 1384 ] = 0; 
		rom[ 1385 ] = 0; 
		rom[ 1386 ] = 0; 
		rom[ 1387 ] = 0; 
		rom[ 1388 ] = 0; 
		rom[ 1389 ] = 8192; 
		rom[ 1390 ] = 8192; 
		rom[ 1391 ] = 0; 
		rom[ 1392 ] = 0; 
		rom[ 1393 ] = 0; 
		rom[ 1394 ] = 0; 
		rom[ 1395 ] = 0; 
		rom[ 1396 ] = 0; 
		rom[ 1397 ] = 0; 
		rom[ 1398 ] = 0; 
		rom[ 1399 ] = 0; 
		rom[ 1400 ] = 0; 
		rom[ 1401 ] = 0; 
		rom[ 1402 ] = 0; 
		rom[ 1403 ] = 0; 
		rom[ 1404 ] = 0; 
		rom[ 1405 ] = 0; 
		rom[ 1406 ] = 0; 
		rom[ 1407 ] = 8192; 
		rom[ 1408 ] = 8192; 
		rom[ 1409 ] = 0; 
		rom[ 1410 ] = 0; 
		rom[ 1411 ] = 8192; 
		rom[ 1412 ] = 0; 
		rom[ 1413 ] = 0; 
		rom[ 1414 ] = 0; 
		rom[ 1415 ] = 0; 
		rom[ 1416 ] = 0; 
		rom[ 1417 ] = 0; 
		rom[ 1418 ] = 0; 
		rom[ 1419 ] = 0; 
		rom[ 1420 ] = 0; 
		rom[ 1421 ] = 0; 
		rom[ 1422 ] = 0; 
		rom[ 1423 ] = 0; 
		rom[ 1424 ] = 8192; 
		rom[ 1425 ] = 0; 
		rom[ 1426 ] = 0; 
		rom[ 1427 ] = 8192; 
		rom[ 1428 ] = 0; 
		rom[ 1429 ] = 0; 
		rom[ 1430 ] = 0; 
		rom[ 1431 ] = 0; 
		rom[ 1432 ] = 0; 
		rom[ 1433 ] = 0; 
		rom[ 1434 ] = 0; 
		rom[ 1435 ] = 0; 
		rom[ 1436 ] = 0; 
		rom[ 1437 ] = 0; 
		rom[ 1438 ] = 0; 
		rom[ 1439 ] = 0; 
		rom[ 1440 ] = 0; 
		rom[ 1441 ] = 0; 
		rom[ 1442 ] = 0; 
		rom[ 1443 ] = 0; 
		rom[ 1444 ] = 0; 
		rom[ 1445 ] = 0; 
		rom[ 1446 ] = 0; 
		rom[ 1447 ] = 0; 
		rom[ 1448 ] = 8192; 
		rom[ 1449 ] = 0; 
		rom[ 1450 ] = 0; 
		rom[ 1451 ] = 8192; 
		rom[ 1452 ] = 0; 
		rom[ 1453 ] = 0; 
		rom[ 1454 ] = 0; 
		rom[ 1455 ] = 0; 
		rom[ 1456 ] = 0; 
		rom[ 1457 ] = 0; 
		rom[ 1458 ] = 0; 
		rom[ 1459 ] = 8192; 
		rom[ 1460 ] = 0; 
		rom[ 1461 ] = 0; 
		rom[ 1462 ] = 0; 
		rom[ 1463 ] = 0; 
		rom[ 1464 ] = 0; 
		rom[ 1465 ] = 0; 
		rom[ 1466 ] = 0; 
		rom[ 1467 ] = 0; 
		rom[ 1468 ] = 8192; 
		rom[ 1469 ] = 8192; 
		rom[ 1470 ] = 8192; 
		rom[ 1471 ] = 0; 
		rom[ 1472 ] = 8192; 
		rom[ 1473 ] = 0; 
		rom[ 1474 ] = 0; 
		rom[ 1475 ] = 0; 
		rom[ 1476 ] = 0; 
		rom[ 1477 ] = 0; 
		rom[ 1478 ] = 0; 
		rom[ 1479 ] = 0; 
		rom[ 1480 ] = 0; 
		rom[ 1481 ] = 0; 
		rom[ 1482 ] = 8192; 
		rom[ 1483 ] = 8192; 
		rom[ 1484 ] = 8192; 
		rom[ 1485 ] = 8192; 
		rom[ 1486 ] = 0; 
		rom[ 1487 ] = 8192; 
		rom[ 1488 ] = 8192; 
		rom[ 1489 ] = 8192; 
		rom[ 1490 ] = 8192; 
		rom[ 1491 ] = 8192; 
		rom[ 1492 ] = 0; 
		rom[ 1493 ] = 8192; 
		rom[ 1494 ] = 0; 
		rom[ 1495 ] = 0; 
		rom[ 1496 ] = 8192; 
		rom[ 1497 ] = 8192; 
		rom[ 1498 ] = 0; 
		rom[ 1499 ] = 0; 
		rom[ 1500 ] = 8192; 
		rom[ 1501 ] = 0; 
		rom[ 1502 ] = 8192; 
		rom[ 1503 ] = 8192; 
		rom[ 1504 ] = 8192; 
		rom[ 1505 ] = 8192; 
		rom[ 1506 ] = 0; 
		rom[ 1507 ] = 0; 
		rom[ 1508 ] = 0; 
		rom[ 1509 ] = 0; 
		rom[ 1510 ] = 8192; 
		rom[ 1511 ] = 8192; 
		rom[ 1512 ] = 0; 
		rom[ 1513 ] = 8192; 
		rom[ 1514 ] = 0; 
		rom[ 1515 ] = 8192; 
		rom[ 1516 ] = 0; 
		rom[ 1517 ] = 0; 
		rom[ 1518 ] = 0; 
		rom[ 1519 ] = 0; 
		rom[ 1520 ] = 8192; 
		rom[ 1521 ] = 8192; 
		rom[ 1522 ] = 0; 
		rom[ 1523 ] = 0; 
		rom[ 1524 ] = 0; 
		rom[ 1525 ] = 0; 
		rom[ 1526 ] = 0; 
		rom[ 1527 ] = 0; 
		rom[ 1528 ] = 0; 
		rom[ 1529 ] = 0; 
		rom[ 1530 ] = 8192; 
		rom[ 1531 ] = 0; 
		rom[ 1532 ] = 0; 
		rom[ 1533 ] = 0; 
		rom[ 1534 ] = 0; 
		rom[ 1535 ] = 0; 
		rom[ 1536 ] = 0; 
		rom[ 1537 ] = 0; 
		rom[ 1538 ] = 0; 
		rom[ 1539 ] = 0; 
		rom[ 1540 ] = 0; 
		rom[ 1541 ] = 0; 
		rom[ 1542 ] = 8192; 
		rom[ 1543 ] = 0; 
		rom[ 1544 ] = 0; 
		rom[ 1545 ] = 0; 
		rom[ 1546 ] = 0; 
		rom[ 1547 ] = 0; 
		rom[ 1548 ] = 8192; 
		rom[ 1549 ] = 0; 
		rom[ 1550 ] = 0; 
		rom[ 1551 ] = 0; 
		rom[ 1552 ] = 0; 
		rom[ 1553 ] = 0; 
		rom[ 1554 ] = 0; 
		rom[ 1555 ] = 0; 
		rom[ 1556 ] = 8192; 
		rom[ 1557 ] = 0; 
		rom[ 1558 ] = 0; 
		rom[ 1559 ] = 0; 
		rom[ 1560 ] = 0; 
		rom[ 1561 ] = 0; 
		rom[ 1562 ] = 0; 
		rom[ 1563 ] = 0; 
		rom[ 1564 ] = 0; 
		rom[ 1565 ] = 8192; 
		rom[ 1566 ] = 8192; 
		rom[ 1567 ] = 0; 
		rom[ 1568 ] = 0; 
		rom[ 1569 ] = 0; 
		rom[ 1570 ] = 0; 
		rom[ 1571 ] = 8192; 
		rom[ 1572 ] = 0; 
		rom[ 1573 ] = 0; 
		rom[ 1574 ] = 0; 
		rom[ 1575 ] = 0; 
		rom[ 1576 ] = 8192; 
		rom[ 1577 ] = 8192; 
		rom[ 1578 ] = 0; 
		rom[ 1579 ] = 0; 
		rom[ 1580 ] = 0; 
		rom[ 1581 ] = 0; 
		rom[ 1582 ] = 0; 
		rom[ 1583 ] = 8192; 
		rom[ 1584 ] = 0; 
		rom[ 1585 ] = 0; 
		rom[ 1586 ] = 0; 
		rom[ 1587 ] = 0; 
		rom[ 1588 ] = 0; 
		rom[ 1589 ] = 0; 
		rom[ 1590 ] = 0; 
		rom[ 1591 ] = 0; 
		rom[ 1592 ] = 0; 
		rom[ 1593 ] = 0; 
		rom[ 1594 ] = 0; 
		rom[ 1595 ] = 0; 
		rom[ 1596 ] = 8192; 
		rom[ 1597 ] = 0; 
		rom[ 1598 ] = 0; 
		rom[ 1599 ] = 0; 
		rom[ 1600 ] = 0; 
		rom[ 1601 ] = 0; 
		rom[ 1602 ] = 0; 
		rom[ 1603 ] = 0; 
		rom[ 1604 ] = 0; 
		rom[ 1605 ] = 8192; 
		rom[ 1606 ] = 0; 
		rom[ 1607 ] = 8192; 
		rom[ 1608 ] = 0; 
		rom[ 1609 ] = 0; 
		rom[ 1610 ] = 8192; 
		rom[ 1611 ] = 0; 
		rom[ 1612 ] = 8192; 
		rom[ 1613 ] = 0; 
		rom[ 1614 ] = 0; 
		rom[ 1615 ] = 0; 
		rom[ 1616 ] = 0; 
		rom[ 1617 ] = 0; 
		rom[ 1618 ] = 0; 
		rom[ 1619 ] = 0; 
		rom[ 1620 ] = 0; 
		rom[ 1621 ] = 0; 
		rom[ 1622 ] = 0; 
		rom[ 1623 ] = 0; 
		rom[ 1624 ] = 0; 
		rom[ 1625 ] = 0; 
		rom[ 1626 ] = 0; 
		rom[ 1627 ] = 0; 
		rom[ 1628 ] = 0; 
		rom[ 1629 ] = 0; 
		rom[ 1630 ] = 0; 
		rom[ 1631 ] = 0; 
		rom[ 1632 ] = 0; 
		rom[ 1633 ] = 0; 
		rom[ 1634 ] = 0; 
		rom[ 1635 ] = 0; 
		rom[ 1636 ] = 0; 
		rom[ 1637 ] = 0; 
		rom[ 1638 ] = 0; 
		rom[ 1639 ] = 0; 
		rom[ 1640 ] = 0; 
		rom[ 1641 ] = 0; 
		rom[ 1642 ] = 0; 
		rom[ 1643 ] = 0; 
		rom[ 1644 ] = 0; 
		rom[ 1645 ] = 0; 
		rom[ 1646 ] = 0; 
		rom[ 1647 ] = 0; 
		rom[ 1648 ] = 8192; 
		rom[ 1649 ] = 0; 
		rom[ 1650 ] = 0; 
		rom[ 1651 ] = 8192; 
		rom[ 1652 ] = 8192; 
		rom[ 1653 ] = 8192; 
		rom[ 1654 ] = 0; 
		rom[ 1655 ] = 0; 
		rom[ 1656 ] = 0; 
		rom[ 1657 ] = 8192; 
		rom[ 1658 ] = 8192; 
		rom[ 1659 ] = 0; 
		rom[ 1660 ] = 8192; 
		rom[ 1661 ] = 0; 
		rom[ 1662 ] = 0; 
		rom[ 1663 ] = 0; 
		rom[ 1664 ] = 0; 
		rom[ 1665 ] = 0; 
		rom[ 1666 ] = 0; 
		rom[ 1667 ] = 0; 
		rom[ 1668 ] = 8192; 
		rom[ 1669 ] = 8192; 
		rom[ 1670 ] = 0; 
		rom[ 1671 ] = 0; 
		rom[ 1672 ] = 0; 
		rom[ 1673 ] = 0; 
		rom[ 1674 ] = 0; 
		rom[ 1675 ] = 0; 
		rom[ 1676 ] = 0; 
		rom[ 1677 ] = 8192; 
		rom[ 1678 ] = 0; 
		rom[ 1679 ] = 0; 
		rom[ 1680 ] = 8192; 
		rom[ 1681 ] = 0; 
		rom[ 1682 ] = 0; 
		rom[ 1683 ] = 8192; 
		rom[ 1684 ] = 8192; 
		rom[ 1685 ] = 8192; 
		rom[ 1686 ] = 0; 
		rom[ 1687 ] = 0; 
		rom[ 1688 ] = 0; 
		rom[ 1689 ] = 0; 
		rom[ 1690 ] = 0; 
		rom[ 1691 ] = 0; 
		rom[ 1692 ] = 0; 
		rom[ 1693 ] = 0; 
		rom[ 1694 ] = 0; 
		rom[ 1695 ] = 0; 
		rom[ 1696 ] = 0; 
		rom[ 1697 ] = 0; 
		rom[ 1698 ] = 0; 
		rom[ 1699 ] = 0; 
		rom[ 1700 ] = 0; 
		rom[ 1701 ] = 0; 
		rom[ 1702 ] = 8192; 
		rom[ 1703 ] = 0; 
		rom[ 1704 ] = 0; 
		rom[ 1705 ] = 0; 
		rom[ 1706 ] = 0; 
		rom[ 1707 ] = 0; 
		rom[ 1708 ] = 0; 
		rom[ 1709 ] = 0; 
		rom[ 1710 ] = 0; 
		rom[ 1711 ] = 0; 
		rom[ 1712 ] = 0; 
		rom[ 1713 ] = 8192; 
		rom[ 1714 ] = 0; 
		rom[ 1715 ] = 0; 
		rom[ 1716 ] = 0; 
		rom[ 1717 ] = 0; 
		rom[ 1718 ] = 0; 
		rom[ 1719 ] = 0; 
		rom[ 1720 ] = 8192; 
		rom[ 1721 ] = 0; 
		rom[ 1722 ] = 0; 
		rom[ 1723 ] = 0; 
		rom[ 1724 ] = 0; 
		rom[ 1725 ] = 0; 
		rom[ 1726 ] = 8192; 
		rom[ 1727 ] = 0; 
		rom[ 1728 ] = 0; 
		rom[ 1729 ] = 0; 
		rom[ 1730 ] = 0; 
		rom[ 1731 ] = 0; 
		rom[ 1732 ] = 0; 
		rom[ 1733 ] = 0; 
		rom[ 1734 ] = 0; 
		rom[ 1735 ] = 0; 
		rom[ 1736 ] = 0; 
		rom[ 1737 ] = 0; 
		rom[ 1738 ] = 0; 
		rom[ 1739 ] = 0; 
		rom[ 1740 ] = 0; 
		rom[ 1741 ] = 0; 
		rom[ 1742 ] = 0; 
		rom[ 1743 ] = 0; 
		rom[ 1744 ] = 0; 
		rom[ 1745 ] = 0; 
		rom[ 1746 ] = 0; 
		rom[ 1747 ] = 0; 
		rom[ 1748 ] = 0; 
		rom[ 1749 ] = 0; 
		rom[ 1750 ] = 0; 
		rom[ 1751 ] = 8192; 
		rom[ 1752 ] = 0; 
		rom[ 1753 ] = 0; 
		rom[ 1754 ] = 0; 
		rom[ 1755 ] = 0; 
		rom[ 1756 ] = 0; 
		rom[ 1757 ] = 0; 
		rom[ 1758 ] = 0; 
		rom[ 1759 ] = 0; 
		rom[ 1760 ] = 0; 
		rom[ 1761 ] = 0; 
		rom[ 1762 ] = 0; 
		rom[ 1763 ] = 8192; 
		rom[ 1764 ] = 8192; 
		rom[ 1765 ] = 0; 
		rom[ 1766 ] = 8192; 
		rom[ 1767 ] = 0; 
		rom[ 1768 ] = 8192; 
		rom[ 1769 ] = 8192; 
		rom[ 1770 ] = 0; 
		rom[ 1771 ] = 0; 
		rom[ 1772 ] = 0; 
		rom[ 1773 ] = 0; 
		rom[ 1774 ] = 0; 
		rom[ 1775 ] = 0; 
		rom[ 1776 ] = 0; 
		rom[ 1777 ] = 0; 
		rom[ 1778 ] = 0; 
		rom[ 1779 ] = 0; 
		rom[ 1780 ] = 0; 
		rom[ 1781 ] = 0; 
		rom[ 1782 ] = 0; 
		rom[ 1783 ] = 0; 
		rom[ 1784 ] = 0; 
		rom[ 1785 ] = 0; 
		rom[ 1786 ] = 8192; 
		rom[ 1787 ] = 0; 
		rom[ 1788 ] = 0; 
		rom[ 1789 ] = 8192; 
		rom[ 1790 ] = 0; 
		rom[ 1791 ] = 8192; 
		rom[ 1792 ] = 0; 
		rom[ 1793 ] = 0; 
		rom[ 1794 ] = 0; 
		rom[ 1795 ] = 0; 
		rom[ 1796 ] = 0; 
		rom[ 1797 ] = 0; 
		rom[ 1798 ] = 0; 
		rom[ 1799 ] = 0; 
		rom[ 1800 ] = 8192; 
		rom[ 1801 ] = 0; 
		rom[ 1802 ] = 0; 
		rom[ 1803 ] = 0; 
		rom[ 1804 ] = 0; 
		rom[ 1805 ] = 8192; 
		rom[ 1806 ] = 0; 
		rom[ 1807 ] = 0; 
		rom[ 1808 ] = 0; 
		rom[ 1809 ] = 0; 
		rom[ 1810 ] = 8192; 
		rom[ 1811 ] = 0; 
		rom[ 1812 ] = 0; 
		rom[ 1813 ] = 8192; 
		rom[ 1814 ] = 0; 
		rom[ 1815 ] = 0; 
		rom[ 1816 ] = 8192; 
		rom[ 1817 ] = 0; 
		rom[ 1818 ] = 0; 
		rom[ 1819 ] = 0; 
		rom[ 1820 ] = 8192; 
		rom[ 1821 ] = 8192; 
		rom[ 1822 ] = 0; 
		rom[ 1823 ] = 0; 
		rom[ 1824 ] = 0; 
		rom[ 1825 ] = 0; 
		rom[ 1826 ] = 0; 
		rom[ 1827 ] = 0; 
		rom[ 1828 ] = 0; 
		rom[ 1829 ] = 0; 
		rom[ 1830 ] = 8192; 
		rom[ 1831 ] = 0; 
		rom[ 1832 ] = 0; 
		rom[ 1833 ] = 8192; 
		rom[ 1834 ] = 0; 
		rom[ 1835 ] = 0; 
		rom[ 1836 ] = 0; 
		rom[ 1837 ] = 8192; 
		rom[ 1838 ] = 8192; 
		rom[ 1839 ] = 0; 
		rom[ 1840 ] = 8192; 
		rom[ 1841 ] = 8192; 
		rom[ 1842 ] = 0; 
		rom[ 1843 ] = 0; 
		rom[ 1844 ] = 0; 
		rom[ 1845 ] = 0; 
		rom[ 1846 ] = 0; 
		rom[ 1847 ] = 0; 
		rom[ 1848 ] = 0; 
		rom[ 1849 ] = 0; 
		rom[ 1850 ] = 0; 
		rom[ 1851 ] = 0; 
		rom[ 1852 ] = 0; 
		rom[ 1853 ] = 0; 
		rom[ 1854 ] = 0; 
		rom[ 1855 ] = 0; 
		rom[ 1856 ] = 0; 
		rom[ 1857 ] = 0; 
		rom[ 1858 ] = 0; 
		rom[ 1859 ] = 0; 
		rom[ 1860 ] = 0; 
		rom[ 1861 ] = 0; 
		rom[ 1862 ] = 8192; 
		rom[ 1863 ] = 0; 
		rom[ 1864 ] = 0; 
		rom[ 1865 ] = 0; 
		rom[ 1866 ] = 0; 
		rom[ 1867 ] = 0; 
		rom[ 1868 ] = 0; 
		rom[ 1869 ] = 0; 
		rom[ 1870 ] = 0; 
		rom[ 1871 ] = 0; 
		rom[ 1872 ] = 0; 
		rom[ 1873 ] = 0; 
		rom[ 1874 ] = 8192; 
		rom[ 1875 ] = 0; 
		rom[ 1876 ] = 0; 
		rom[ 1877 ] = 0; 
		rom[ 1878 ] = 0; 
		rom[ 1879 ] = 0; 
		rom[ 1880 ] = 8192; 
		rom[ 1881 ] = 0; 
		rom[ 1882 ] = 0; 
		rom[ 1883 ] = 8192; 
		rom[ 1884 ] = 8192; 
		rom[ 1885 ] = 0; 
		rom[ 1886 ] = 0; 
		rom[ 1887 ] = 0; 
		rom[ 1888 ] = 0; 
		rom[ 1889 ] = 0; 
		rom[ 1890 ] = 0; 
		rom[ 1891 ] = 0; 
		rom[ 1892 ] = 8192; 
		rom[ 1893 ] = 8192; 
		rom[ 1894 ] = 0; 
		rom[ 1895 ] = 0; 
		rom[ 1896 ] = 0; 
		rom[ 1897 ] = 0; 
		rom[ 1898 ] = 0; 
		rom[ 1899 ] = 0; 
		rom[ 1900 ] = 8192; 
		rom[ 1901 ] = 8192; 
		rom[ 1902 ] = 0; 
		rom[ 1903 ] = 0; 
		rom[ 1904 ] = 0; 
		rom[ 1905 ] = 0; 
		rom[ 1906 ] = 0; 
		rom[ 1907 ] = 0; 
		rom[ 1908 ] = 0; 
		rom[ 1909 ] = 0; 
		rom[ 1910 ] = 0; 
		rom[ 1911 ] = 0; 
		rom[ 1912 ] = 0; 
		rom[ 1913 ] = 8192; 
		rom[ 1914 ] = 8192; 
		rom[ 1915 ] = 8192; 
		rom[ 1916 ] = 0; 
		rom[ 1917 ] = 8192; 
		rom[ 1918 ] = 0; 
		rom[ 1919 ] = 0; 
		rom[ 1920 ] = 0; 
		rom[ 1921 ] = 0; 
		rom[ 1922 ] = 0; 
		rom[ 1923 ] = 0; 
		rom[ 1924 ] = 0; 
		rom[ 1925 ] = 0; 
		rom[ 1926 ] = 0; 
		rom[ 1927 ] = 0; 
		rom[ 1928 ] = 0; 
		rom[ 1929 ] = 0; 
		rom[ 1930 ] = 0; 
		rom[ 1931 ] = 0; 
		rom[ 1932 ] = 0; 
		rom[ 1933 ] = 0; 
		rom[ 1934 ] = 0; 
		rom[ 1935 ] = 0; 
		rom[ 1936 ] = 0; 
		rom[ 1937 ] = 0; 
		rom[ 1938 ] = 0; 
		rom[ 1939 ] = 0; 
		rom[ 1940 ] = 8192; 
		rom[ 1941 ] = 0; 
		rom[ 1942 ] = 0; 
		rom[ 1943 ] = 0; 
		rom[ 1944 ] = 0; 
		rom[ 1945 ] = 0; 
		rom[ 1946 ] = 8192; 
		rom[ 1947 ] = 8192; 
		rom[ 1948 ] = 0; 
		rom[ 1949 ] = 8192; 
		rom[ 1950 ] = 8192; 
		rom[ 1951 ] = 8192; 
		rom[ 1952 ] = 0; 
		rom[ 1953 ] = 0; 
		rom[ 1954 ] = 0; 
		rom[ 1955 ] = 0; 
		rom[ 1956 ] = 8192; 
		rom[ 1957 ] = 0; 
		rom[ 1958 ] = 8192; 
		rom[ 1959 ] = 0; 
		rom[ 1960 ] = 0; 
		rom[ 1961 ] = 0; 
		rom[ 1962 ] = 0; 
		rom[ 1963 ] = 8192; 
		rom[ 1964 ] = 0; 
		rom[ 1965 ] = 0; 
		rom[ 1966 ] = 0; 
		rom[ 1967 ] = 8192; 
		rom[ 1968 ] = 0; 
		rom[ 1969 ] = 0; 
		rom[ 1970 ] = 0; 
		rom[ 1971 ] = 0; 
		rom[ 1972 ] = 0; 
		rom[ 1973 ] = 0; 
		rom[ 1974 ] = 0; 
		rom[ 1975 ] = 0; 
		rom[ 1976 ] = 0; 
		rom[ 1977 ] = 0; 
		rom[ 1978 ] = 8192; 
		rom[ 1979 ] = 0; 
		rom[ 1980 ] = 0; 
		rom[ 1981 ] = 0; 
		rom[ 1982 ] = 0; 
		rom[ 1983 ] = 0; 
		rom[ 1984 ] = 0; 
		rom[ 1985 ] = 8192; 
		rom[ 1986 ] = 0; 
		rom[ 1987 ] = 0; 
		rom[ 1988 ] = 0; 
		rom[ 1989 ] = 0; 
		rom[ 1990 ] = 0; 
		rom[ 1991 ] = 0; 
		rom[ 1992 ] = 8192; 
		rom[ 1993 ] = 0; 
		rom[ 1994 ] = 0; 
		rom[ 1995 ] = 0; 
		rom[ 1996 ] = 0; 
		rom[ 1997 ] = 0; 
		rom[ 1998 ] = 0; 
		rom[ 1999 ] = 0; 
		rom[ 2000 ] = 0; 
		rom[ 2001 ] = 0; 
		rom[ 2002 ] = 0; 
		rom[ 2003 ] = 8192; 
		rom[ 2004 ] = 8192; 
		rom[ 2005 ] = 8192; 
		rom[ 2006 ] = 0; 
		rom[ 2007 ] = 0; 
		rom[ 2008 ] = 0; 
		rom[ 2009 ] = 8192; 
		rom[ 2010 ] = 0; 
		rom[ 2011 ] = 0; 
		rom[ 2012 ] = 0; 
		rom[ 2013 ] = 0; 
		rom[ 2014 ] = 0; 
		rom[ 2015 ] = 8192; 
		rom[ 2016 ] = 0; 
		rom[ 2017 ] = 8192; 
		rom[ 2018 ] = 0; 
		rom[ 2019 ] = 8192; 
		rom[ 2020 ] = 8192; 
		rom[ 2021 ] = 8192; 
		rom[ 2022 ] = 0; 
		rom[ 2023 ] = 0; 
		rom[ 2024 ] = 0; 
		rom[ 2025 ] = 8192; 
		rom[ 2026 ] = 0; 
		rom[ 2027 ] = 0; 
		rom[ 2028 ] = 0; 
		rom[ 2029 ] = 0; 
		rom[ 2030 ] = 0; 
		rom[ 2031 ] = 0; 
		rom[ 2032 ] = 0; 
		rom[ 2033 ] = 0; 
		rom[ 2034 ] = 0; 
		rom[ 2035 ] = 0; 
		rom[ 2036 ] = 8192; 
		rom[ 2037 ] = 0; 
		rom[ 2038 ] = 0; 
		rom[ 2039 ] = 8192; 
		rom[ 2040 ] = 8192; 
		rom[ 2041 ] = 8192; 
		rom[ 2042 ] = 8192; 
		rom[ 2043 ] = 0; 
		rom[ 2044 ] = 0; 
		rom[ 2045 ] = 0; 
		rom[ 2046 ] = 8192; 
		rom[ 2047 ] = 8192; 
		rom[ 2048 ] = 0; 
		rom[ 2049 ] = 0; 
		rom[ 2050 ] = 0; 
		rom[ 2051 ] = 0; 
		rom[ 2052 ] = 0; 
		rom[ 2053 ] = 0; 
		rom[ 2054 ] = 0; 
		rom[ 2055 ] = 0; 
		rom[ 2056 ] = 0; 
		rom[ 2057 ] = 0; 
		rom[ 2058 ] = 0; 
		rom[ 2059 ] = 0; 
		rom[ 2060 ] = 0; 
		rom[ 2061 ] = 8192; 
		rom[ 2062 ] = 0; 
		rom[ 2063 ] = 0; 
		rom[ 2064 ] = 0; 
		rom[ 2065 ] = 0; 
		rom[ 2066 ] = 0; 
		rom[ 2067 ] = 8192; 
		rom[ 2068 ] = 0; 
		rom[ 2069 ] = 0; 
		rom[ 2070 ] = 8192; 
		rom[ 2071 ] = 0; 
		rom[ 2072 ] = 8192; 
		rom[ 2073 ] = 8192; 
		rom[ 2074 ] = 8192; 
		rom[ 2075 ] = 0; 
		rom[ 2076 ] = 8192; 
		rom[ 2077 ] = 0; 
		rom[ 2078 ] = 0; 
		rom[ 2079 ] = 0; 
		rom[ 2080 ] = 0; 
		rom[ 2081 ] = 0; 
		rom[ 2082 ] = 0; 
		rom[ 2083 ] = 0; 
		rom[ 2084 ] = 8192; 
		rom[ 2085 ] = 0; 
		rom[ 2086 ] = 0; 
		rom[ 2087 ] = 0; 
		rom[ 2088 ] = 0; 
		rom[ 2089 ] = 8192; 
		rom[ 2090 ] = 8192; 
		rom[ 2091 ] = 8192; 
		rom[ 2092 ] = 8192; 
		rom[ 2093 ] = 0; 
		rom[ 2094 ] = 0; 
		rom[ 2095 ] = 8192; 
		rom[ 2096 ] = 8192; 
		rom[ 2097 ] = 0; 
		rom[ 2098 ] = 0; 
		rom[ 2099 ] = 0; 
		rom[ 2100 ] = 0; 
		rom[ 2101 ] = 0; 
		rom[ 2102 ] = 8192; 
		rom[ 2103 ] = 8192; 
		rom[ 2104 ] = 8192; 
		rom[ 2105 ] = 8192; 
		rom[ 2106 ] = 8192; 
		rom[ 2107 ] = 0; 
		rom[ 2108 ] = 0; 
		rom[ 2109 ] = 0; 
		rom[ 2110 ] = 0; 
		rom[ 2111 ] = 0; 
		rom[ 2112 ] = 0; 
		rom[ 2113 ] = 0; 
		rom[ 2114 ] = 0; 
		rom[ 2115 ] = 0; 
		rom[ 2116 ] = 0; 
		rom[ 2117 ] = 0; 
		rom[ 2118 ] = 0; 
		rom[ 2119 ] = 0; 
		rom[ 2120 ] = 0; 
		rom[ 2121 ] = 0; 
		rom[ 2122 ] = 0; 
		rom[ 2123 ] = 0; 
		rom[ 2124 ] = 0; 
		rom[ 2125 ] = 0; 
		rom[ 2126 ] = 0; 
		rom[ 2127 ] = 0; 
		rom[ 2128 ] = 0; 
		rom[ 2129 ] = 0; 
		rom[ 2130 ] = 0; 
		rom[ 2131 ] = 0; 
		rom[ 2132 ] = 0; 
		rom[ 2133 ] = 0; 
		rom[ 2134 ] = 0; 
		rom[ 2135 ] = 0; 
		rom[ 2136 ] = 0; 
		rom[ 2137 ] = 0; 
		rom[ 2138 ] = 0; 
		rom[ 2139 ] = 0; 
		rom[ 2140 ] = 0; 
		rom[ 2141 ] = 0; 
		rom[ 2142 ] = 8192; 
		rom[ 2143 ] = 0; 
		rom[ 2144 ] = 0; 
		rom[ 2145 ] = 0; 
		rom[ 2146 ] = 8192; 
		rom[ 2147 ] = 0; 
		rom[ 2148 ] = 0; 
		rom[ 2149 ] = 0; 
		rom[ 2150 ] = 0; 
		rom[ 2151 ] = 0; 
		rom[ 2152 ] = 0; 
		rom[ 2153 ] = 8192; 
		rom[ 2154 ] = 0; 
		rom[ 2155 ] = 0; 
		rom[ 2156 ] = 0; 
		rom[ 2157 ] = 0; 
		rom[ 2158 ] = 0; 
		rom[ 2159 ] = 0; 
		rom[ 2160 ] = 0; 
		rom[ 2161 ] = 0; 
		rom[ 2162 ] = 0; 
		rom[ 2163 ] = 0; 
		rom[ 2164 ] = 8192; 
		rom[ 2165 ] = 8192; 
		rom[ 2166 ] = 8192; 
		rom[ 2167 ] = 8192; 
		rom[ 2168 ] = 0; 
		rom[ 2169 ] = 0; 
		rom[ 2170 ] = 8192; 
		rom[ 2171 ] = 0; 
		rom[ 2172 ] = 0; 
		rom[ 2173 ] = 0; 
		rom[ 2174 ] = 8192; 
		rom[ 2175 ] = 0; 
		rom[ 2176 ] = 0; 
		rom[ 2177 ] = 0; 
		rom[ 2178 ] = 0; 
		rom[ 2179 ] = 0; 
		rom[ 2180 ] = 0; 
		rom[ 2181 ] = 8192; 
		rom[ 2182 ] = 0; 
		rom[ 2183 ] = 0; 
		rom[ 2184 ] = 0; 
		rom[ 2185 ] = 0; 
		rom[ 2186 ] = 8192; 
		rom[ 2187 ] = 0; 
		rom[ 2188 ] = 0; 
		rom[ 2189 ] = 8192; 
		rom[ 2190 ] = 0; 
		rom[ 2191 ] = 0; 
		rom[ 2192 ] = 8192; 
		rom[ 2193 ] = 0; 
		rom[ 2194 ] = 0; 
		rom[ 2195 ] = 0; 
		rom[ 2196 ] = 0; 
		rom[ 2197 ] = 8192; 
		rom[ 2198 ] = 0; 
		rom[ 2199 ] = 8192; 
		rom[ 2200 ] = 0; 
		rom[ 2201 ] = 0; 
		rom[ 2202 ] = 0; 
		rom[ 2203 ] = 0; 
		rom[ 2204 ] = 8192; 
		rom[ 2205 ] = 8192; 
		rom[ 2206 ] = 8192; 
		rom[ 2207 ] = 0; 
		rom[ 2208 ] = 0; 
		rom[ 2209 ] = 0; 
		rom[ 2210 ] = 0; 
		rom[ 2211 ] = 0; 
		rom[ 2212 ] = 0; 
		rom[ 2213 ] = 0; 
		rom[ 2214 ] = 0; 
		rom[ 2215 ] = 0; 
		rom[ 2216 ] = 0; 
		rom[ 2217 ] = 0; 
		rom[ 2218 ] = 0; 
		rom[ 2219 ] = 0; 
		rom[ 2220 ] = 0; 
		rom[ 2221 ] = 0; 
		rom[ 2222 ] = 0; 
		rom[ 2223 ] = 0; 
		rom[ 2224 ] = 0; 
		rom[ 2225 ] = 0; 
		rom[ 2226 ] = 0; 
		rom[ 2227 ] = 0; 
		rom[ 2228 ] = 0; 
		rom[ 2229 ] = 0; 
		rom[ 2230 ] = 8192; 
		rom[ 2231 ] = 0; 
		rom[ 2232 ] = 0; 
		rom[ 2233 ] = 0; 
		rom[ 2234 ] = 0; 
		rom[ 2235 ] = 0; 
		rom[ 2236 ] = 0; 
		rom[ 2237 ] = 0; 
		rom[ 2238 ] = 8192; 
		rom[ 2239 ] = 0; 
		rom[ 2240 ] = 0; 
		rom[ 2241 ] = 0; 
		rom[ 2242 ] = 0; 
		rom[ 2243 ] = 0; 
		rom[ 2244 ] = 0; 
		rom[ 2245 ] = 8192; 
		rom[ 2246 ] = 0; 
		rom[ 2247 ] = 0; 
		rom[ 2248 ] = 0; 
		rom[ 2249 ] = 0; 
		rom[ 2250 ] = 0; 
		rom[ 2251 ] = 0; 
		rom[ 2252 ] = 8192; 
		rom[ 2253 ] = 8192; 
		rom[ 2254 ] = 0; 
		rom[ 2255 ] = 0; 
		rom[ 2256 ] = 0; 
		rom[ 2257 ] = 0; 
		rom[ 2258 ] = 0; 
		rom[ 2259 ] = 0; 
		rom[ 2260 ] = 0; 
		rom[ 2261 ] = 0; 
		rom[ 2262 ] = 0; 
		rom[ 2263 ] = 0; 
		rom[ 2264 ] = 8192; 
		rom[ 2265 ] = 8192; 
		rom[ 2266 ] = 0; 
		rom[ 2267 ] = 0; 
		rom[ 2268 ] = 0; 
		rom[ 2269 ] = 0; 
		rom[ 2270 ] = 0; 
		rom[ 2271 ] = 0; 
		rom[ 2272 ] = 0; 
		rom[ 2273 ] = 8192; 
		rom[ 2274 ] = 0; 
		rom[ 2275 ] = 8192; 
		rom[ 2276 ] = 0; 
		rom[ 2277 ] = 0; 
		rom[ 2278 ] = 8192; 
		rom[ 2279 ] = 8192; 
		rom[ 2280 ] = 0; 
		rom[ 2281 ] = 0; 
		rom[ 2282 ] = 0; 
		rom[ 2283 ] = 0; 
		rom[ 2284 ] = 0; 
		rom[ 2285 ] = 0; 
		rom[ 2286 ] = 0; 
		rom[ 2287 ] = 8192; 
		rom[ 2288 ] = 0; 
		rom[ 2289 ] = 8192; 
		rom[ 2290 ] = 8192; 
		rom[ 2291 ] = 8192; 
		rom[ 2292 ] = 8192; 
		rom[ 2293 ] = 0; 
		rom[ 2294 ] = 0; 
		rom[ 2295 ] = 0; 
		rom[ 2296 ] = 0; 
		rom[ 2297 ] = 0; 
		rom[ 2298 ] = 0; 
		rom[ 2299 ] = 0; 
		rom[ 2300 ] = 0; 
		rom[ 2301 ] = 0; 
		rom[ 2302 ] = 0; 
		rom[ 2303 ] = 0; 
		rom[ 2304 ] = 0; 
		rom[ 2305 ] = 0; 
		rom[ 2306 ] = 0; 
		rom[ 2307 ] = 0; 
		rom[ 2308 ] = 0; 
		rom[ 2309 ] = 0; 
		rom[ 2310 ] = 0; 
		rom[ 2311 ] = 0; 
		rom[ 2312 ] = 0; 
		rom[ 2313 ] = 0; 
		rom[ 2314 ] = 0; 
		rom[ 2315 ] = 0; 
		rom[ 2316 ] = 0; 
		rom[ 2317 ] = 0; 
		rom[ 2318 ] = 8192; 
		rom[ 2319 ] = 0; 
		rom[ 2320 ] = 8192; 
		rom[ 2321 ] = 8192; 
		rom[ 2322 ] = 8192; 
		rom[ 2323 ] = 0; 
		rom[ 2324 ] = 0; 
		rom[ 2325 ] = 0; 
		rom[ 2326 ] = 0; 
		rom[ 2327 ] = 0; 
		rom[ 2328 ] = 0; 
		rom[ 2329 ] = 8192; 
		rom[ 2330 ] = 0; 
		rom[ 2331 ] = 0; 
		rom[ 2332 ] = 0; 
		rom[ 2333 ] = 0; 
		rom[ 2334 ] = 0; 
		rom[ 2335 ] = 0; 
		rom[ 2336 ] = 0; 
		rom[ 2337 ] = 8192; 
		rom[ 2338 ] = 8192; 
		rom[ 2339 ] = 8192; 
		rom[ 2340 ] = 0; 
		rom[ 2341 ] = 8192; 
		rom[ 2342 ] = 0; 
		rom[ 2343 ] = 0; 
		rom[ 2344 ] = 0; 
		rom[ 2345 ] = 0; 
		rom[ 2346 ] = 8192; 
		rom[ 2347 ] = 8192; 
		rom[ 2348 ] = 0; 
		rom[ 2349 ] = 0; 
		rom[ 2350 ] = 8192; 
		rom[ 2351 ] = 8192; 
		rom[ 2352 ] = 0; 
		rom[ 2353 ] = 0; 
		rom[ 2354 ] = 8192; 
		rom[ 2355 ] = 0; 
		rom[ 2356 ] = 8192; 
		rom[ 2357 ] = 0; 
		rom[ 2358 ] = 0; 
		rom[ 2359 ] = 0; 
		rom[ 2360 ] = 0; 
		rom[ 2361 ] = 0; 
		rom[ 2362 ] = 0; 
		rom[ 2363 ] = 0; 
		rom[ 2364 ] = 0; 
		rom[ 2365 ] = 8192; 
		rom[ 2366 ] = 0; 
		rom[ 2367 ] = 0; 
		rom[ 2368 ] = 8192; 
		rom[ 2369 ] = 8192; 
		rom[ 2370 ] = 0; 
		rom[ 2371 ] = 0; 
		rom[ 2372 ] = 0; 
		rom[ 2373 ] = 0; 
		rom[ 2374 ] = 8192; 
		rom[ 2375 ] = 0; 
		rom[ 2376 ] = 0; 
		rom[ 2377 ] = 0; 
		rom[ 2378 ] = 8192; 
		rom[ 2379 ] = 0; 
		rom[ 2380 ] = 0; 
		rom[ 2381 ] = 0; 
		rom[ 2382 ] = 8192; 
		rom[ 2383 ] = 8192; 
		rom[ 2384 ] = 0; 
		rom[ 2385 ] = 0; 
		rom[ 2386 ] = 8192; 
		rom[ 2387 ] = 0; 
		rom[ 2388 ] = 0; 
		rom[ 2389 ] = 0; 
		rom[ 2390 ] = 0; 
		rom[ 2391 ] = 0; 
		rom[ 2392 ] = 0; 
		rom[ 2393 ] = 0; 
		rom[ 2394 ] = 0; 
		rom[ 2395 ] = 8192; 
		rom[ 2396 ] = 0; 
		rom[ 2397 ] = 0; 
		rom[ 2398 ] = 0; 
		rom[ 2399 ] = 0; 
		rom[ 2400 ] = 0; 
		rom[ 2401 ] = 0; 
		rom[ 2402 ] = 0; 
		rom[ 2403 ] = 0; 
		rom[ 2404 ] = 0; 
		rom[ 2405 ] = 0; 
		rom[ 2406 ] = 0; 
		rom[ 2407 ] = 0; 
		rom[ 2408 ] = 0; 
		rom[ 2409 ] = 0; 
		rom[ 2410 ] = 0; 
		rom[ 2411 ] = 0; 
		rom[ 2412 ] = 8192; 
		rom[ 2413 ] = 0; 
		rom[ 2414 ] = 0; 
		rom[ 2415 ] = 0; 
		rom[ 2416 ] = 0; 
		rom[ 2417 ] = 0; 
		rom[ 2418 ] = 0; 
		rom[ 2419 ] = 0; 
		rom[ 2420 ] = 0; 
		rom[ 2421 ] = 0; 
		rom[ 2422 ] = 0; 
		rom[ 2423 ] = 0; 
		rom[ 2424 ] = 0; 
		rom[ 2425 ] = 8192; 
		rom[ 2426 ] = 0; 
		rom[ 2427 ] = 0; 
		rom[ 2428 ] = 8192; 
		rom[ 2429 ] = 8192; 
		rom[ 2430 ] = 0; 
		rom[ 2431 ] = 0; 
		rom[ 2432 ] = 0; 
		rom[ 2433 ] = 8192; 
		rom[ 2434 ] = 0; 
		rom[ 2435 ] = 0; 
		rom[ 2436 ] = 8192; 
		rom[ 2437 ] = 8192; 
		rom[ 2438 ] = 8192; 
		rom[ 2439 ] = 0; 
		rom[ 2440 ] = 0; 
		rom[ 2441 ] = 8192; 
		rom[ 2442 ] = 0; 
		rom[ 2443 ] = 0; 
		rom[ 2444 ] = 0; 
		rom[ 2445 ] = 8192; 
		rom[ 2446 ] = 0; 
		rom[ 2447 ] = 0; 
		rom[ 2448 ] = 8192; 
		rom[ 2449 ] = 0; 
		rom[ 2450 ] = 0; 
		rom[ 2451 ] = 0; 
		rom[ 2452 ] = 0; 
		rom[ 2453 ] = 0; 
		rom[ 2454 ] = 0; 
		rom[ 2455 ] = 0; 
		rom[ 2456 ] = 8192; 
		rom[ 2457 ] = 8192; 
		rom[ 2458 ] = 0; 
		rom[ 2459 ] = 0; 
		rom[ 2460 ] = 8192; 
		rom[ 2461 ] = 0; 
		rom[ 2462 ] = 0; 
		rom[ 2463 ] = 8192; 
		rom[ 2464 ] = 0; 
		rom[ 2465 ] = 0; 
		rom[ 2466 ] = 0; 
		rom[ 2467 ] = 0; 
		rom[ 2468 ] = 0; 
		rom[ 2469 ] = 0; 
		rom[ 2470 ] = 0; 
		rom[ 2471 ] = 0; 
		rom[ 2472 ] = 0; 
		rom[ 2473 ] = 0; 
		rom[ 2474 ] = 0; 
		rom[ 2475 ] = 0; 
		rom[ 2476 ] = 0; 
		rom[ 2477 ] = 0; 
		rom[ 2478 ] = 0; 
		rom[ 2479 ] = 8192; 
		rom[ 2480 ] = 0; 
		rom[ 2481 ] = 0; 
		rom[ 2482 ] = 0; 
		rom[ 2483 ] = 0; 
		rom[ 2484 ] = 0; 
		rom[ 2485 ] = 8192; 
		rom[ 2486 ] = 0; 
		rom[ 2487 ] = 0; 
		rom[ 2488 ] = 0; 
		rom[ 2489 ] = 0; 
		rom[ 2490 ] = 8192; 
		rom[ 2491 ] = 8192; 
		rom[ 2492 ] = 8192; 
		rom[ 2493 ] = 8192; 
		rom[ 2494 ] = 0; 
		rom[ 2495 ] = 0; 
		rom[ 2496 ] = 8192; 
		rom[ 2497 ] = 0; 
		rom[ 2498 ] = 0; 
		rom[ 2499 ] = 0; 
		rom[ 2500 ] = 0; 
		rom[ 2501 ] = 8192; 
		rom[ 2502 ] = 0; 
		rom[ 2503 ] = 0; 
		rom[ 2504 ] = 0; 
		rom[ 2505 ] = 0; 
		rom[ 2506 ] = 0; 
		rom[ 2507 ] = 0; 
		rom[ 2508 ] = 0; 
		rom[ 2509 ] = 0; 
		rom[ 2510 ] = 8192; 
		rom[ 2511 ] = 8192; 
		rom[ 2512 ] = 0; 
		rom[ 2513 ] = 8192; 
		rom[ 2514 ] = 0; 
		rom[ 2515 ] = 0; 
		rom[ 2516 ] = 0; 
		rom[ 2517 ] = 0; 
		rom[ 2518 ] = 0; 
		rom[ 2519 ] = 0; 
		rom[ 2520 ] = 0; 
		rom[ 2521 ] = 0; 
		rom[ 2522 ] = 0; 
		rom[ 2523 ] = 0; 
		rom[ 2524 ] = 0; 
		rom[ 2525 ] = 0; 
		rom[ 2526 ] = 0; 
		rom[ 2527 ] = 0; 
		rom[ 2528 ] = 0; 
		rom[ 2529 ] = 0; 
		rom[ 2530 ] = 0; 
		rom[ 2531 ] = 0; 
		rom[ 2532 ] = 0; 
		rom[ 2533 ] = 0; 
		rom[ 2534 ] = 0; 
		rom[ 2535 ] = 8192; 
		rom[ 2536 ] = 8192; 
		rom[ 2537 ] = 8192; 
		rom[ 2538 ] = 0; 
		rom[ 2539 ] = 8192; 
		rom[ 2540 ] = 8192; 
		rom[ 2541 ] = 0; 
		rom[ 2542 ] = 8192; 
		rom[ 2543 ] = 8192; 
		rom[ 2544 ] = 8192; 
		rom[ 2545 ] = 0; 
		rom[ 2546 ] = 0; 
		rom[ 2547 ] = 0; 
		rom[ 2548 ] = 0; 
		rom[ 2549 ] = 0; 
		rom[ 2550 ] = 0; 
		rom[ 2551 ] = 0; 
		rom[ 2552 ] = 0; 
		rom[ 2553 ] = 8192; 
		rom[ 2554 ] = 0; 
		rom[ 2555 ] = 8192; 
		rom[ 2556 ] = 0; 
		rom[ 2557 ] = 0; 
		rom[ 2558 ] = 0; 
		rom[ 2559 ] = 0; 
		rom[ 2560 ] = 0; 
		rom[ 2561 ] = 0; 
		rom[ 2562 ] = 0; 
		rom[ 2563 ] = 0; 
		rom[ 2564 ] = 0; 
		rom[ 2565 ] = 0; 
		rom[ 2566 ] = 0; 
		rom[ 2567 ] = 0; 
		rom[ 2568 ] = 8192; 
		rom[ 2569 ] = 0; 
		rom[ 2570 ] = 0; 
		rom[ 2571 ] = 0; 
		rom[ 2572 ] = 0; 
		rom[ 2573 ] = 0; 
		rom[ 2574 ] = 0; 
		rom[ 2575 ] = 0; 
		rom[ 2576 ] = 0; 
		rom[ 2577 ] = 0; 
		rom[ 2578 ] = 0; 
		rom[ 2579 ] = 0; 
		rom[ 2580 ] = 8192; 
		rom[ 2581 ] = 8192; 
		rom[ 2582 ] = 8192; 
		rom[ 2583 ] = 8192; 
		rom[ 2584 ] = 8192; 
		rom[ 2585 ] = 0; 
		rom[ 2586 ] = 0; 
		rom[ 2587 ] = 8192; 
		rom[ 2588 ] = 0; 
		rom[ 2589 ] = 8192; 
		rom[ 2590 ] = 8192; 
		rom[ 2591 ] = 0; 
		rom[ 2592 ] = 8192; 
		rom[ 2593 ] = 0; 
		rom[ 2594 ] = 0; 
		rom[ 2595 ] = 8192; 
		rom[ 2596 ] = 0; 
		rom[ 2597 ] = 8192; 
		rom[ 2598 ] = 8192; 
		rom[ 2599 ] = 0; 
		rom[ 2600 ] = 0; 
		rom[ 2601 ] = 0; 
		rom[ 2602 ] = 0; 
		rom[ 2603 ] = 0; 
		rom[ 2604 ] = 0; 
		rom[ 2605 ] = 0; 
		rom[ 2606 ] = 0; 
		rom[ 2607 ] = 0; 
		rom[ 2608 ] = 8192; 
		rom[ 2609 ] = 0; 
		rom[ 2610 ] = 0; 
		rom[ 2611 ] = 8192; 
		rom[ 2612 ] = 8192; 
		rom[ 2613 ] = 0; 
		rom[ 2614 ] = 0; 
		rom[ 2615 ] = 0; 
		rom[ 2616 ] = 8192; 
		rom[ 2617 ] = 0; 
		rom[ 2618 ] = 0; 
		rom[ 2619 ] = 0; 
		rom[ 2620 ] = 0; 
		rom[ 2621 ] = 0; 
		rom[ 2622 ] = 0; 
		rom[ 2623 ] = 0; 
		rom[ 2624 ] = 0; 
		rom[ 2625 ] = 0; 
		rom[ 2626 ] = 8192; 
		rom[ 2627 ] = 0; 
		rom[ 2628 ] = 0; 
		rom[ 2629 ] = 0; 
		rom[ 2630 ] = 0; 
		rom[ 2631 ] = 0; 
		rom[ 2632 ] = 0; 
		rom[ 2633 ] = 0; 
		rom[ 2634 ] = 0; 
		rom[ 2635 ] = 0; 
		rom[ 2636 ] = 0; 
		rom[ 2637 ] = 0; 
		rom[ 2638 ] = 0; 
		rom[ 2639 ] = 0; 
		rom[ 2640 ] = 0; 
		rom[ 2641 ] = 8192; 
		rom[ 2642 ] = 8192; 
		rom[ 2643 ] = 0; 
		rom[ 2644 ] = 0; 
		rom[ 2645 ] = 8192; 
		rom[ 2646 ] = 8192; 
		rom[ 2647 ] = 0; 
		rom[ 2648 ] = 8192; 
		rom[ 2649 ] = 0; 
		rom[ 2650 ] = 0; 
		rom[ 2651 ] = 0; 
		rom[ 2652 ] = 0; 
		rom[ 2653 ] = 8192; 
		rom[ 2654 ] = 0; 
		rom[ 2655 ] = 0; 
		rom[ 2656 ] = 8192; 
		rom[ 2657 ] = 0; 
		rom[ 2658 ] = 0; 
		rom[ 2659 ] = 0; 
		rom[ 2660 ] = 0; 
		rom[ 2661 ] = 0; 
		rom[ 2662 ] = 0; 
		rom[ 2663 ] = 0; 
		rom[ 2664 ] = 0; 
		rom[ 2665 ] = 0; 
		rom[ 2666 ] = 0; 
		rom[ 2667 ] = 0; 
		rom[ 2668 ] = 0; 
		rom[ 2669 ] = 0; 
		rom[ 2670 ] = 8192; 
		rom[ 2671 ] = 8192; 
		rom[ 2672 ] = 0; 
		rom[ 2673 ] = 0; 
		rom[ 2674 ] = 8192; 
		rom[ 2675 ] = 8192; 
		rom[ 2676 ] = 0; 
		rom[ 2677 ] = 0; 
		rom[ 2678 ] = 0; 
		rom[ 2679 ] = 8192; 
		rom[ 2680 ] = 0; 
		rom[ 2681 ] = 0; 
		rom[ 2682 ] = 0; 
		rom[ 2683 ] = 0; 
		rom[ 2684 ] = 0; 
		rom[ 2685 ] = 0; 
		rom[ 2686 ] = 0; 
		rom[ 2687 ] = 0; 
		rom[ 2688 ] = 0; 
		rom[ 2689 ] = 0; 
		rom[ 2690 ] = 0; 
		rom[ 2691 ] = 0; 
		rom[ 2692 ] = 0; 
		rom[ 2693 ] = 0; 
		rom[ 2694 ] = 0; 
		rom[ 2695 ] = 0; 
		rom[ 2696 ] = 0; 
		rom[ 2697 ] = 0; 
		rom[ 2698 ] = 0; 
		rom[ 2699 ] = 0; 
		rom[ 2700 ] = 0; 
		rom[ 2701 ] = 0; 
		rom[ 2702 ] = 0; 
		rom[ 2703 ] = 0; 
		rom[ 2704 ] = 0; 
		rom[ 2705 ] = 0; 
		rom[ 2706 ] = 8192; 
		rom[ 2707 ] = 8192; 
		rom[ 2708 ] = 0; 
		rom[ 2709 ] = 0; 
		rom[ 2710 ] = 0; 
		rom[ 2711 ] = 8192; 
		rom[ 2712 ] = 0; 
		rom[ 2713 ] = 0; 
		rom[ 2714 ] = 0; 
		rom[ 2715 ] = 0; 
		rom[ 2716 ] = 0; 
		rom[ 2717 ] = 0; 
		rom[ 2718 ] = 8192; 
		rom[ 2719 ] = 0; 
		rom[ 2720 ] = 0; 
		rom[ 2721 ] = 0; 
		rom[ 2722 ] = 0; 
		rom[ 2723 ] = 8192; 
		rom[ 2724 ] = 0; 
		rom[ 2725 ] = 0; 
		rom[ 2726 ] = 0; 
		rom[ 2727 ] = 0; 
		rom[ 2728 ] = 8192; 
		rom[ 2729 ] = 0; 
		rom[ 2730 ] = 0; 
		rom[ 2731 ] = 0; 
		rom[ 2732 ] = 0; 
		rom[ 2733 ] = 0; 
		rom[ 2734 ] = 0; 
		rom[ 2735 ] = 0; 
		rom[ 2736 ] = 0; 
		rom[ 2737 ] = 0; 
		rom[ 2738 ] = 0; 
		rom[ 2739 ] = 0; 
		rom[ 2740 ] = 0; 
		rom[ 2741 ] = 0; 
		rom[ 2742 ] = 0; 
		rom[ 2743 ] = 0; 
		rom[ 2744 ] = 0; 
		rom[ 2745 ] = 0; 
		rom[ 2746 ] = 0; 
		rom[ 2747 ] = 0; 
		rom[ 2748 ] = 0; 
		rom[ 2749 ] = 0; 
		rom[ 2750 ] = 0; 
		rom[ 2751 ] = 0; 
		rom[ 2752 ] = 0; 
		rom[ 2753 ] = 0; 
		rom[ 2754 ] = 0; 
		rom[ 2755 ] = 0; 
		rom[ 2756 ] = 0; 
		rom[ 2757 ] = 8192; 
		rom[ 2758 ] = 0; 
		rom[ 2759 ] = 8192; 
		rom[ 2760 ] = 0; 
		rom[ 2761 ] = 0; 
		rom[ 2762 ] = 0; 
		rom[ 2763 ] = 0; 
		rom[ 2764 ] = 0; 
		rom[ 2765 ] = 0; 
		rom[ 2766 ] = 0; 
		rom[ 2767 ] = 0; 
		rom[ 2768 ] = 0; 
		rom[ 2769 ] = 8192; 
		rom[ 2770 ] = 8192; 
		rom[ 2771 ] = 8192; 
		rom[ 2772 ] = 0; 
		rom[ 2773 ] = 0; 
		rom[ 2774 ] = 8192; 
		rom[ 2775 ] = 0; 
		rom[ 2776 ] = 8192; 
		rom[ 2777 ] = 8192; 
		rom[ 2778 ] = 8192; 
		rom[ 2779 ] = 8192; 
		rom[ 2780 ] = 0; 
		rom[ 2781 ] = 0; 
		rom[ 2782 ] = 0; 
		rom[ 2783 ] = 0; 
		rom[ 2784 ] = 0; 
		rom[ 2785 ] = 0; 
		rom[ 2786 ] = 8192; 
		rom[ 2787 ] = 0; 
		rom[ 2788 ] = 0; 
		rom[ 2789 ] = 0; 
		rom[ 2790 ] = 0; 
		rom[ 2791 ] = 0; 
		rom[ 2792 ] = 0; 
		rom[ 2793 ] = 0; 
		rom[ 2794 ] = 8192; 
		rom[ 2795 ] = 8192; 
		rom[ 2796 ] = 0; 
		rom[ 2797 ] = 8192; 
		rom[ 2798 ] = 8192; 
		rom[ 2799 ] = 8192; 
		rom[ 2800 ] = 8192; 
		rom[ 2801 ] = 8192; 
		rom[ 2802 ] = 0; 
		rom[ 2803 ] = 0; 
		rom[ 2804 ] = 0; 
		rom[ 2805 ] = 0; 
		rom[ 2806 ] = 0; 
		rom[ 2807 ] = 0; 
		rom[ 2808 ] = 0; 
		rom[ 2809 ] = 0; 
		rom[ 2810 ] = 0; 
		rom[ 2811 ] = 0; 
		rom[ 2812 ] = 0; 
		rom[ 2813 ] = 0; 
		rom[ 2814 ] = 0; 
		rom[ 2815 ] = 0; 
		rom[ 2816 ] = 8192; 
		rom[ 2817 ] = 8192; 
		rom[ 2818 ] = 0; 
		rom[ 2819 ] = 0; 
		rom[ 2820 ] = 0; 
		rom[ 2821 ] = 0; 
		rom[ 2822 ] = 0; 
		rom[ 2823 ] = 0; 
		rom[ 2824 ] = 0; 
		rom[ 2825 ] = 0; 
		rom[ 2826 ] = 8192; 
		rom[ 2827 ] = 0; 
		rom[ 2828 ] = 0; 
		rom[ 2829 ] = 0; 
		rom[ 2830 ] = 0; 
		rom[ 2831 ] = 0; 
		rom[ 2832 ] = 8192; 
		rom[ 2833 ] = 0; 
		rom[ 2834 ] = 0; 
		rom[ 2835 ] = 0; 
		rom[ 2836 ] = 0; 
		rom[ 2837 ] = 0; 
		rom[ 2838 ] = 8192; 
		rom[ 2839 ] = 0; 
		rom[ 2840 ] = 0; 
		rom[ 2841 ] = 0; 
		rom[ 2842 ] = 0; 
		rom[ 2843 ] = 0; 
		rom[ 2844 ] = 0; 
		rom[ 2845 ] = 0; 
		rom[ 2846 ] = 8192; 
		rom[ 2847 ] = 0; 
		rom[ 2848 ] = 0; 
		rom[ 2849 ] = 0; 
		rom[ 2850 ] = 0; 
		rom[ 2851 ] = 8192; 
		rom[ 2852 ] = 0; 
		rom[ 2853 ] = 0; 
		rom[ 2854 ] = 0; 
		rom[ 2855 ] = 0; 
		rom[ 2856 ] = 0; 
		rom[ 2857 ] = 8192; 
		rom[ 2858 ] = 8192; 
		rom[ 2859 ] = 0; 
		rom[ 2860 ] = 0; 
		rom[ 2861 ] = 0; 
		rom[ 2862 ] = 0; 
		rom[ 2863 ] = 0; 
		rom[ 2864 ] = 0; 
		rom[ 2865 ] = 0; 
		rom[ 2866 ] = 8192; 
		rom[ 2867 ] = 0; 
		rom[ 2868 ] = 0; 
		rom[ 2869 ] = 0; 
		rom[ 2870 ] = 0; 
		rom[ 2871 ] = 0; 
		rom[ 2872 ] = 0; 
		rom[ 2873 ] = 0; 
		rom[ 2874 ] = 0; 
		rom[ 2875 ] = 8192; 
		rom[ 2876 ] = 8192; 
		rom[ 2877 ] = 8192; 
		rom[ 2878 ] = 8192; 
		rom[ 2879 ] = 8192; 
		rom[ 2880 ] = 8192; 
		rom[ 2881 ] = 8192; 
		rom[ 2882 ] = 8192; 
		rom[ 2883 ] = 8192; 
		rom[ 2884 ] = 0; 
		rom[ 2885 ] = 0; 
		rom[ 2886 ] = 0; 
		rom[ 2887 ] = 0; 
		rom[ 2888 ] = 0; 
		rom[ 2889 ] = 0; 
		rom[ 2890 ] = 0; 
		rom[ 2891 ] = 0; 
		rom[ 2892 ] = 0; 
		rom[ 2893 ] = 0; 
		rom[ 2894 ] = 8192; 
		rom[ 2895 ] = 8192; 
		rom[ 2896 ] = 0; 
		rom[ 2897 ] = 0; 
		rom[ 2898 ] = 8192; 
		rom[ 2899 ] = 8192; 
		rom[ 2900 ] = 0; 
		rom[ 2901 ] = 8192; 
		rom[ 2902 ] = 0; 
		rom[ 2903 ] = 0; 
		rom[ 2904 ] = 0; 
		rom[ 2905 ] = 0; 
		rom[ 2906 ] = 0; 
		rom[ 2907 ] = 0; 
		rom[ 2908 ] = 0; 
		rom[ 2909 ] = 0; 
		rom[ 2910 ] = 0; 
		rom[ 2911 ] = 0; 
		rom[ 2912 ] = 8192; 
	
	end
endmodule

module weak_thresh_rom(
	input 				clk,
	input		[11:0]	addr,
	output reg	[12:0]	q    // x y w h 5bit*4
	);
	reg					[12:0]	rom [4095:0];
	always @(posedge clk) q <= rom[addr];
	initial begin
		rom[ 0    ] =   -129;
		rom[ 1    ] =     50;
		rom[ 2    ] =     89;
		rom[ 3    ] =     23;
		rom[ 4    ] =     61;
		rom[ 5    ] =    407;
		rom[ 6    ] =     11;
		rom[ 7    ] =    -77;
		rom[ 8    ] =     24;
		rom[ 9    ] =    -86;
		rom[ 10   ] =     83;
		rom[ 11   ] =     87;
		rom[ 12   ] =    375;
		rom[ 13   ] =    148;
		rom[ 14   ] =    -78;
		rom[ 15   ] =     33;
		rom[ 16   ] =     75;
		rom[ 17   ] =    -28;
		rom[ 18   ] =    -40;
		rom[ 19   ] =     64;
		rom[ 20   ] =    -84;
		rom[ 21   ] =   -563;
		rom[ 22   ] =     58;
		rom[ 23   ] =     41;
		rom[ 24   ] =    374;
		rom[ 25   ] =    285;
		rom[ 26   ] =    129;
		rom[ 27   ] =     58;
		rom[ 28   ] =     59;
		rom[ 29   ] =    -12;
		rom[ 30   ] =    134;
		rom[ 31   ] =    -29;
		rom[ 32   ] =    206;
		rom[ 33   ] =    192;
		rom[ 34   ] =   -284;
		rom[ 35   ] =   -200;
		rom[ 36   ] =    347;
		rom[ 37   ] =     -7;
		rom[ 38   ] =    473;
		rom[ 39   ] =   -210;
		rom[ 40   ] =   -174;
		rom[ 41   ] =   1522;
		rom[ 42   ] =     79;
		rom[ 43   ] =     71;
		rom[ 44   ] =    162;
		rom[ 45   ] =    -37;
		rom[ 46   ] =      7;
		rom[ 47   ] =    123;
		rom[ 48   ] =   -322;
		rom[ 49   ] =      8;
		rom[ 50   ] =    110;
		rom[ 51   ] =   -184;
		rom[ 52   ] =   -269;
		rom[ 53   ] =     64;
		rom[ 54   ] =    596;
		rom[ 55   ] =     25;
		rom[ 56   ] =     27;
		rom[ 57   ] =     75;
		rom[ 58   ] =     81;
		rom[ 59   ] =  -1136;
		rom[ 60   ] =     37;
		rom[ 61   ] =   -154;
		rom[ 62   ] =     75;
		rom[ 63   ] =    -45;
		rom[ 64   ] =    138;
		rom[ 65   ] =   -146;
		rom[ 66   ] =    -46;
		rom[ 67   ] =   -267;
		rom[ 68   ] =   -173;
		rom[ 69   ] =      7;
		rom[ 70   ] =   -529;
		rom[ 71   ] =     93;
		rom[ 72   ] =   -139;
		rom[ 73   ] =    107;
		rom[ 74   ] =     91;
		rom[ 75   ] =    -23;
		rom[ 76   ] =    178;
		rom[ 77   ] =    234;
		rom[ 78   ] =      9;
		rom[ 79   ] =     53;
		rom[ 80   ] =   -108;
		rom[ 81   ] =    -23;
		rom[ 82   ] =    -67;
		rom[ 83   ] =   -279;
		rom[ 84   ] =    163;
		rom[ 85   ] =    770;
		rom[ 86   ] =    319;
		rom[ 87   ] =      0;
		rom[ 88   ] =    348;
		rom[ 89   ] =     36;
		rom[ 90   ] =     36;
		rom[ 91   ] =    -96;
		rom[ 92   ] =     28;
		rom[ 93   ] =    138;
		rom[ 94   ] =    -13;
		rom[ 95   ] =    119;
		rom[ 96   ] =    -34;
		rom[ 97   ] =    -44;
		rom[ 98   ] =   -100;
		rom[ 99   ] =     15;
		rom[ 100  ] =    -50;
		rom[ 101  ] =    -19;
		rom[ 102  ] =    314;
		rom[ 103  ] =    117;
		rom[ 104  ] =     80;
		rom[ 105  ] =   -119;
		rom[ 106  ] =   -119;
		rom[ 107  ] =     80;
		rom[ 108  ] =     17;
		rom[ 109  ] =   -145;
		rom[ 110  ] =    -66;
		rom[ 111  ] =    -90;
		rom[ 112  ] =    -93;
		rom[ 113  ] =     68;
		rom[ 114  ] =    -54;
		rom[ 115  ] =   -138;
		rom[ 116  ] =     69;
		rom[ 117  ] =     13;
		rom[ 118  ] =    342;
		rom[ 119  ] =   1056;
		rom[ 120  ] =   -149;
		rom[ 121  ] =    -67;
		rom[ 122  ] =    -15;
		rom[ 123  ] =    -26;
		rom[ 124  ] =    -15;
		rom[ 125  ] =   -186;
		rom[ 126  ] =    -98;
		rom[ 127  ] =   -317;
		rom[ 128  ] =     96;
		rom[ 129  ] =    -10;
		rom[ 130  ] =    491;
		rom[ 131  ] =      9;
		rom[ 132  ] =    285;
		rom[ 133  ] =   -191;
		rom[ 134  ] =   -205;
		rom[ 135  ] =    123;
		rom[ 136  ] =    373;
		rom[ 137  ] =     52;
		rom[ 138  ] =     65;
		rom[ 139  ] =      9;
		rom[ 140  ] =    130;
		rom[ 141  ] =     11;
		rom[ 142  ] =    -49;
		rom[ 143  ] =     87;
		rom[ 144  ] =    124;
		rom[ 145  ] =   -184;
		rom[ 146  ] =   -293;
		rom[ 147  ] =    242;
		rom[ 148  ] =     27;
		rom[ 149  ] =    168;
		rom[ 150  ] =     -3;
		rom[ 151  ] =   -124;
		rom[ 152  ] =    -52;
		rom[ 153  ] =    153;
		rom[ 154  ] =    100;
		rom[ 155  ] =    233;
		rom[ 156  ] =    -66;
		rom[ 157  ] =   -722;
		rom[ 158  ] =    721;
		rom[ 159  ] =    -30;
		rom[ 160  ] =    249;
		rom[ 161  ] =   -119;
		rom[ 162  ] =   -186;
		rom[ 163  ] =    152;
		rom[ 164  ] =    -99;
		rom[ 165  ] =   -244;
		rom[ 166  ] =   -123;
		rom[ 167  ] =     30;
		rom[ 168  ] =     -8;
		rom[ 169  ] =     85;
		rom[ 170  ] =    -27;
		rom[ 171  ] =     76;
		rom[ 172  ] =   -181;
		rom[ 173  ] =     93;
		rom[ 174  ] =     -4;
		rom[ 175  ] =     70;
		rom[ 176  ] =   -141;
		rom[ 177  ] =    274;
		rom[ 178  ] =    973;
		rom[ 179  ] =    -52;
		rom[ 180  ] =     43;
		rom[ 181  ] =     69;
		rom[ 182  ] =    -29;
		rom[ 183  ] =     43;
		rom[ 184  ] =     25;
		rom[ 185  ] =     53;
		rom[ 186  ] =     12;
		rom[ 187  ] =   -447;
		rom[ 188  ] =     33;
		rom[ 189  ] =    128;
		rom[ 190  ] =    130;
		rom[ 191  ] =     27;
		rom[ 192  ] =    107;
		rom[ 193  ] =     52;
		rom[ 194  ] =    107;
		rom[ 195  ] =    -61;
		rom[ 196  ] =   -159;
		rom[ 197  ] =    -23;
		rom[ 198  ] =     -6;
		rom[ 199  ] =   -116;
		rom[ 200  ] =    271;
		rom[ 201  ] =     36;
		rom[ 202  ] =     46;
		rom[ 203  ] =    -11;
		rom[ 204  ] =     46;
		rom[ 205  ] =     29;
		rom[ 206  ] =    130;
		rom[ 207  ] =    103;
		rom[ 208  ] =     30;
		rom[ 209  ] =    134;
		rom[ 210  ] =    -11;
		rom[ 211  ] =   -155;
		rom[ 212  ] =   -159;
		rom[ 213  ] =     11;
		rom[ 214  ] =   -221;
		rom[ 215  ] =    -34;
		rom[ 216  ] =    138;
		rom[ 217  ] =   -460;
		rom[ 218  ] =    -42;
		rom[ 219  ] =    -20;
		rom[ 220  ] =    -38;
		rom[ 221  ] =    -48;
		rom[ 222  ] =    -95;
		rom[ 223  ] =     69;
		rom[ 224  ] =    -98;
		rom[ 225  ] =   -151;
		rom[ 226  ] =   -252;
		rom[ 227  ] =     88;
		rom[ 228  ] =    -15;
		rom[ 229  ] =    183;
		rom[ 230  ] =    234;
		rom[ 231  ] =    -46;
		rom[ 232  ] =    -49;
		rom[ 233  ] =     92;
		rom[ 234  ] =    -81;
		rom[ 235  ] =     65;
		rom[ 236  ] =    -37;
		rom[ 237  ] =    -18;
		rom[ 238  ] =    521;
		rom[ 239  ] =    195;
		rom[ 240  ] =    219;
		rom[ 241  ] =   -162;
		rom[ 242  ] =   -275;
		rom[ 243  ] =    546;
		rom[ 244  ] =   -856;
		rom[ 245  ] =   -268;
		rom[ 246  ] =    253;
		rom[ 247  ] =   -104;
		rom[ 248  ] =   -142;
		rom[ 249  ] =    -74;
		rom[ 250  ] =     61;
		rom[ 251  ] =    189;
		rom[ 252  ] =     63;
		rom[ 253  ] =     52;
		rom[ 254  ] =    201;
		rom[ 255  ] =     51;
		rom[ 256  ] =    -76;
		rom[ 257  ] =    171;
		rom[ 258  ] =   -210;
		rom[ 259  ] =   -290;
		rom[ 260  ] =     68;
		rom[ 261  ] =    -25;
		rom[ 262  ] =   -161;
		rom[ 263  ] =      0;
		rom[ 264  ] =    -91;
		rom[ 265  ] =      7;
		rom[ 266  ] =      4;
		rom[ 267  ] =    160;
		rom[ 268  ] =    254;
		rom[ 269  ] =      8;
		rom[ 270  ] =      3;
		rom[ 271  ] =    -28;
		rom[ 272  ] =    -97;
		rom[ 273  ] =   -420;
		rom[ 274  ] =    -39;
		rom[ 275  ] =    163;
		rom[ 276  ] =    -53;
		rom[ 277  ] =   -207;
		rom[ 278  ] =    102;
		rom[ 279  ] =    -31;
		rom[ 280  ] =    175;
		rom[ 281  ] =      0;
		rom[ 282  ] =     37;
		rom[ 283  ] =     45;
		rom[ 284  ] =   -214;
		rom[ 285  ] =   -942;
		rom[ 286  ] =    -67;
		rom[ 287  ] =    -70;
		rom[ 288  ] =   -150;
		rom[ 289  ] =    -42;
		rom[ 290  ] =    -56;
		rom[ 291  ] =    120;
		rom[ 292  ] =     98;
		rom[ 293  ] =     25;
		rom[ 294  ] =    -91;
		rom[ 295  ] =    -28;
		rom[ 296  ] =   -166;
		rom[ 297  ] =   -100;
		rom[ 298  ] =     10;
		rom[ 299  ] =    -80;
		rom[ 300  ] =   -121;
		rom[ 301  ] =    -61;
		rom[ 302  ] =   -248;
		rom[ 303  ] =    -52;
		rom[ 304  ] =    -82;
		rom[ 305  ] =   -125;
		rom[ 306  ] =    -84;
		rom[ 307  ] =     -7;
		rom[ 308  ] =   -128;
		rom[ 309  ] =     77;
		rom[ 310  ] =     25;
		rom[ 311  ] =    -41;
		rom[ 312  ] =     -5;
		rom[ 313  ] =    -16;
		rom[ 314  ] =   -180;
		rom[ 315  ] =   -248;
		rom[ 316  ] =   -134;
		rom[ 317  ] =   -603;
		rom[ 318  ] =    -48;
		rom[ 319  ] =    594;
		rom[ 320  ] =    210;
		rom[ 321  ] =     12;
		rom[ 322  ] =   -178;
		rom[ 323  ] =    528;
		rom[ 324  ] =   -373;
		rom[ 325  ] =     58;
		rom[ 326  ] =    134;
		rom[ 327  ] =     51;
		rom[ 328  ] =     60;
		rom[ 329  ] =   -137;
		rom[ 330  ] =    583;
		rom[ 331  ] =    -25;
		rom[ 332  ] =     74;
		rom[ 333  ] =    102;
		rom[ 334  ] =    190;
		rom[ 335  ] =    -36;
		rom[ 336  ] =    167;
		rom[ 337  ] =   -140;
		rom[ 338  ] =   -162;
		rom[ 339  ] =     10;
		rom[ 340  ] =    112;
		rom[ 341  ] =    143;
		rom[ 342  ] =     18;
		rom[ 343  ] =     11;
		rom[ 344  ] =    144;
		rom[ 345  ] =    106;
		rom[ 346  ] =    -64;
		rom[ 347  ] =    -31;
		rom[ 348  ] =     85;
		rom[ 349  ] =    245;
		rom[ 350  ] =    159;
		rom[ 351  ] =     88;
		rom[ 352  ] =   -112;
		rom[ 353  ] =     42;
		rom[ 354  ] =    101;
		rom[ 355  ] =    -65;
		rom[ 356  ] =    199;
		rom[ 357  ] =      5;
		rom[ 358  ] =   -360;
		rom[ 359  ] =     75;
		rom[ 360  ] =    144;
		rom[ 361  ] =   -835;
		rom[ 362  ] =    -68;
		rom[ 363  ] =    154;
		rom[ 364  ] =      9;
		rom[ 365  ] =    -60;
		rom[ 366  ] =   -197;
		rom[ 367  ] =   -120;
		rom[ 368  ] =   -189;
		rom[ 369  ] =   -114;
		rom[ 370  ] =    -23;
		rom[ 371  ] =    -41;
		rom[ 372  ] =     46;
		rom[ 373  ] =    212;
		rom[ 374  ] =    136;
		rom[ 375  ] =    -59;
		rom[ 376  ] =   -140;
		rom[ 377  ] =   -330;
		rom[ 378  ] =     -3;
		rom[ 379  ] =    397;
		rom[ 380  ] =    149;
		rom[ 381  ] =    211;
		rom[ 382  ] =   -100;
		rom[ 383  ] =   1340;
		rom[ 384  ] =     31;
		rom[ 385  ] =    662;
		rom[ 386  ] =    -19;
		rom[ 387  ] =    -75;
		rom[ 388  ] =    318;
		rom[ 389  ] =     77;
		rom[ 390  ] =   -325;
		rom[ 391  ] =   -278;
		rom[ 392  ] =    -24;
		rom[ 393  ] =    130;
		rom[ 394  ] =   -122;
		rom[ 395  ] =   -329;
		rom[ 396  ] =     15;
		rom[ 397  ] =    137;
		rom[ 398  ] =     33;
		rom[ 399  ] =    413;
		rom[ 400  ] =    -40;
		rom[ 401  ] =     29;
		rom[ 402  ] =    102;
		rom[ 403  ] =   1143;
		rom[ 404  ] =   -181;
		rom[ 405  ] =    -57;
		rom[ 406  ] =    564;
		rom[ 407  ] =    141;
		rom[ 408  ] =     76;
		rom[ 409  ] =    102;
		rom[ 410  ] =    234;
		rom[ 411  ] =     61;
		rom[ 412  ] =     36;
		rom[ 413  ] =    124;
		rom[ 414  ] =   -180;
		rom[ 415  ] =     75;
		rom[ 416  ] =     43;
		rom[ 417  ] =   -188;
		rom[ 418  ] =    339;
		rom[ 419  ] =    -36;
		rom[ 420  ] =    175;
		rom[ 421  ] =    -35;
		rom[ 422  ] =    -17;
		rom[ 423  ] =     33;
		rom[ 424  ] =    396;
		rom[ 425  ] =   -125;
		rom[ 426  ] =   -249;
		rom[ 427  ] =   -156;
		rom[ 428  ] =    -39;
		rom[ 429  ] =    200;
		rom[ 430  ] =   -170;
		rom[ 431  ] =    -82;
		rom[ 432  ] =     -4;
		rom[ 433  ] =   -137;
		rom[ 434  ] =     79;
		rom[ 435  ] =     -1;
		rom[ 436  ] =     -1;
		rom[ 437  ] =   -382;
		rom[ 438  ] =   -318;
		rom[ 439  ] =     69;
		rom[ 440  ] =    -87;
		rom[ 441  ] =    -52;
		rom[ 442  ] =     32;
		rom[ 443  ] =    421;
		rom[ 444  ] =   -153;
		rom[ 445  ] =    104;
		rom[ 446  ] =      2;
		rom[ 447  ] =  -1182;
		rom[ 448  ] =    373;
		rom[ 449  ] =    493;
		rom[ 450  ] =   -302;
		rom[ 451  ] =   -135;
		rom[ 452  ] =   -179;
		rom[ 453  ] =    741;
		rom[ 454  ] =    -48;
		rom[ 455  ] =     18;
		rom[ 456  ] =     28;
		rom[ 457  ] =    -97;
		rom[ 458  ] =   -275;
		rom[ 459  ] =   -267;
		rom[ 460  ] =     93;
		rom[ 461  ] =    -77;
		rom[ 462  ] =    -28;
		rom[ 463  ] =   -164;
		rom[ 464  ] =   -166;
		rom[ 465  ] =    -50;
		rom[ 466  ] =   -111;
		rom[ 467  ] =   -361;
		rom[ 468  ] =    -32;
		rom[ 469  ] =   -171;
		rom[ 470  ] =    187;
		rom[ 471  ] =   -577;
		rom[ 472  ] =   -242;
		rom[ 473  ] =     17;
		rom[ 474  ] =     -8;
		rom[ 475  ] =   1127;
		rom[ 476  ] =   -108;
		rom[ 477  ] =    167;
		rom[ 478  ] =     22;
		rom[ 479  ] =    130;
		rom[ 480  ] =   -169;
		rom[ 481  ] =   -393;
		rom[ 482  ] =    -47;
		rom[ 483  ] =     75;
		rom[ 484  ] =   -139;
		rom[ 485  ] =   -100;
		rom[ 486  ] =    200;
		rom[ 487  ] =    -84;
		rom[ 488  ] =    -94;
		rom[ 489  ] =    264;
		rom[ 490  ] =     51;
		rom[ 491  ] =    -49;
		rom[ 492  ] =   -108;
		rom[ 493  ] =   -104;
		rom[ 494  ] =    160;
		rom[ 495  ] =    -24;
		rom[ 496  ] =   -139;
		rom[ 497  ] =    166;
		rom[ 498  ] =    104;
		rom[ 499  ] =    817;
		rom[ 500  ] =     50;
		rom[ 501  ] =    160;
		rom[ 502  ] =   -126;
		rom[ 503  ] =   -145;
		rom[ 504  ] =   -252;
		rom[ 505  ] =    -48;
		rom[ 506  ] =    274;
		rom[ 507  ] =    -84;
		rom[ 508  ] =    -91;
		rom[ 509  ] =      4;
		rom[ 510  ] =    146;
		rom[ 511  ] =    125;
		rom[ 512  ] =     22;
		rom[ 513  ] =    -25;
		rom[ 514  ] =   -124;
		rom[ 515  ] =    -39;
		rom[ 516  ] =   -233;
		rom[ 517  ] =     16;
		rom[ 518  ] =    138;
		rom[ 519  ] =   -141;
		rom[ 520  ] =    192;
		rom[ 521  ] =    -35;
		rom[ 522  ] =    268;
		rom[ 523  ] =   -180;
		rom[ 524  ] =     70;
		rom[ 525  ] =    135;
		rom[ 526  ] =    -86;
		rom[ 527  ] =    121;
		rom[ 528  ] =    226;
		rom[ 529  ] =   -137;
		rom[ 530  ] =     80;
		rom[ 531  ] =    -85;
		rom[ 532  ] =    133;
		rom[ 533  ] =    -44;
		rom[ 534  ] =    -40;
		rom[ 535  ] =    -15;
		rom[ 536  ] =   -171;
		rom[ 537  ] =   -140;
		rom[ 538  ] =     41;
		rom[ 539  ] =   -368;
		rom[ 540  ] =    106;
		rom[ 541  ] =    -15;
		rom[ 542  ] =    130;
		rom[ 543  ] =     79;
		rom[ 544  ] =      7;
		rom[ 545  ] =   -180;
		rom[ 546  ] =   -183;
		rom[ 547  ] =   -440;
		rom[ 548  ] =   -526;
		rom[ 549  ] =   -183;
		rom[ 550  ] =   -180;
		rom[ 551  ] =   -502;
		rom[ 552  ] =    -81;
		rom[ 553  ] =    -63;
		rom[ 554  ] =   -200;
		rom[ 555  ] =    229;
		rom[ 556  ] =    -40;
		rom[ 557  ] =     55;
		rom[ 558  ] =     26;
		rom[ 559  ] =     29;
		rom[ 560  ] =     19;
		rom[ 561  ] =     39;
		rom[ 562  ] =   -112;
		rom[ 563  ] =   -161;
		rom[ 564  ] =   -125;
		rom[ 565  ] =     -6;
		rom[ 566  ] =    781;
		rom[ 567  ] =     21;
		rom[ 568  ] =     98;
		rom[ 569  ] =   -108;
		rom[ 570  ] =     22;
		rom[ 571  ] =    222;
		rom[ 572  ] =      0;
		rom[ 573  ] =     62;
		rom[ 574  ] =     69;
		rom[ 575  ] =    124;
		rom[ 576  ] =     26;
		rom[ 577  ] =    580;
		rom[ 578  ] =     79;
		rom[ 579  ] =    -70;
		rom[ 580  ] =    -25;
		rom[ 581  ] =    -65;
		rom[ 582  ] =   -414;
		rom[ 583  ] =    -30;
		rom[ 584  ] =    181;
		rom[ 585  ] =   -476;
		rom[ 586  ] =     19;
		rom[ 587  ] =     91;
		rom[ 588  ] =    -49;
		rom[ 589  ] =    229;
		rom[ 590  ] =    -35;
		rom[ 591  ] =     27;
		rom[ 592  ] =    -74;
		rom[ 593  ] =    -93;
		rom[ 594  ] =     52;
		rom[ 595  ] =    -56;
		rom[ 596  ] =    128;
		rom[ 597  ] =    381;
		rom[ 598  ] =    106;
		rom[ 599  ] =     67;
		rom[ 600  ] =     -7;
		rom[ 601  ] =    -36;
		rom[ 602  ] =     92;
		rom[ 603  ] =   -154;
		rom[ 604  ] =    -22;
		rom[ 605  ] =    -97;
		rom[ 606  ] =   -108;
		rom[ 607  ] =     50;
		rom[ 608  ] =    395;
		rom[ 609  ] =   -112;
		rom[ 610  ] =    -64;
		rom[ 611  ] =     -8;
		rom[ 612  ] =     49;
		rom[ 613  ] =    -63;
		rom[ 614  ] =    -17;
		rom[ 615  ] =    -86;
		rom[ 616  ] =    -69;
		rom[ 617  ] =   -167;
		rom[ 618  ] =    -33;
		rom[ 619  ] =    -78;
		rom[ 620  ] =   -181;
		rom[ 621  ] =   -255;
		rom[ 622  ] =     -4;
		rom[ 623  ] =     97;
		rom[ 624  ] =     87;
		rom[ 625  ] =     82;
		rom[ 626  ] =   -117;
		rom[ 627  ] =     14;
		rom[ 628  ] =    233;
		rom[ 629  ] =   -384;
		rom[ 630  ] =     72;
		rom[ 631  ] =    935;
		rom[ 632  ] =   -749;
		rom[ 633  ] =   -286;
		rom[ 634  ] =     62;
		rom[ 635  ] =     27;
		rom[ 636  ] =    -65;
		rom[ 637  ] =     53;
		rom[ 638  ] =     53;
		rom[ 639  ] =   -163;
		rom[ 640  ] =     61;
		rom[ 641  ] =    -84;
		rom[ 642  ] =    -91;
		rom[ 643  ] =    -32;
		rom[ 644  ] =     62;
		rom[ 645  ] =   -129;
		rom[ 646  ] =   -126;
		rom[ 647  ] =    -63;
		rom[ 648  ] =    144;
		rom[ 649  ] =    -73;
		rom[ 650  ] =    -13;
		rom[ 651  ] =     64;
		rom[ 652  ] =    122;
		rom[ 653  ] =     12;
		rom[ 654  ] =    347;
		rom[ 655  ] =   -240;
		rom[ 656  ] =    183;
		rom[ 657  ] =    165;
		rom[ 658  ] =    154;
		rom[ 659  ] =    248;
		rom[ 660  ] =    -81;
		rom[ 661  ] =   -679;
		rom[ 662  ] =    282;
		rom[ 663  ] =     46;
		rom[ 664  ] =      6;
		rom[ 665  ] =    326;
		rom[ 666  ] =   -234;
		rom[ 667  ] =     30;
		rom[ 668  ] =    -73;
		rom[ 669  ] =    387;
		rom[ 670  ] =     22;
		rom[ 671  ] =     28;
		rom[ 672  ] =    141;
		rom[ 673  ] =   -212;
		rom[ 674  ] =   -283;
		rom[ 675  ] =    -22;
		rom[ 676  ] =    280;
		rom[ 677  ] =   -274;
		rom[ 678  ] =    -86;
		rom[ 679  ] =     83;
		rom[ 680  ] =   -192;
		rom[ 681  ] =    768;
		rom[ 682  ] =   -177;
		rom[ 683  ] =     81;
		rom[ 684  ] =     33;
		rom[ 685  ] =    111;
		rom[ 686  ] =   -375;
		rom[ 687  ] =    -51;
		rom[ 688  ] =     60;
		rom[ 689  ] =    119;
		rom[ 690  ] =     35;
		rom[ 691  ] =   -224;
		rom[ 692  ] =    -60;
		rom[ 693  ] =    102;
		rom[ 694  ] =    190;
		rom[ 695  ] =     72;
		rom[ 696  ] =    668;
		rom[ 697  ] =     53;
		rom[ 698  ] =    -64;
		rom[ 699  ] =    329;
		rom[ 700  ] =    144;
		rom[ 701  ] =    135;
		rom[ 702  ] =     49;
		rom[ 703  ] =    176;
		rom[ 704  ] =    124;
		rom[ 705  ] =    145;
		rom[ 706  ] =    -59;
		rom[ 707  ] =     51;
		rom[ 708  ] =     41;
		rom[ 709  ] =    118;
		rom[ 710  ] =      2;
		rom[ 711  ] =    198;
		rom[ 712  ] =    132;
		rom[ 713  ] =    136;
		rom[ 714  ] =     26;
		rom[ 715  ] =    -23;
		rom[ 716  ] =     52;
		rom[ 717  ] =     24;
		rom[ 718  ] =     10;
		rom[ 719  ] =    -69;
		rom[ 720  ] =    115;
		rom[ 721  ] =     42;
		rom[ 722  ] =     40;
		rom[ 723  ] =    106;
		rom[ 724  ] =   -104;
		rom[ 725  ] =    -14;
		rom[ 726  ] =     37;
		rom[ 727  ] =     86;
		rom[ 728  ] =   -209;
		rom[ 729  ] =   -255;
		rom[ 730  ] =   -135;
		rom[ 731  ] =   -153;
		rom[ 732  ] =    508;
		rom[ 733  ] =    -36;
		rom[ 734  ] =   -245;
		rom[ 735  ] =     25;
		rom[ 736  ] =    -72;
		rom[ 737  ] =     72;
		rom[ 738  ] =     21;
		rom[ 739  ] =    -43;
		rom[ 740  ] =    855;
		rom[ 741  ] =   -108;
		rom[ 742  ] =    241;
		rom[ 743  ] =    -47;
		rom[ 744  ] =    188;
		rom[ 745  ] =    -93;
		rom[ 746  ] =    -33;
		rom[ 747  ] =     14;
		rom[ 748  ] =    202;
		rom[ 749  ] =     14;
		rom[ 750  ] =   -126;
		rom[ 751  ] =    354;
		rom[ 752  ] =   -559;
		rom[ 753  ] =    -23;
		rom[ 754  ] =    -73;
		rom[ 755  ] =    -81;
		rom[ 756  ] =   -235;
		rom[ 757  ] =   -340;
		rom[ 758  ] =   -220;
		rom[ 759  ] =    -34;
		rom[ 760  ] =    226;
		rom[ 761  ] =   -275;
		rom[ 762  ] =    -97;
		rom[ 763  ] =     22;
		rom[ 764  ] =     87;
		rom[ 765  ] =   -100;
		rom[ 766  ] =    -80;
		rom[ 767  ] =   -218;
		rom[ 768  ] =     29;
		rom[ 769  ] =    -92;
		rom[ 770  ] =   -337;
		rom[ 771  ] =    536;
		rom[ 772  ] =     58;
		rom[ 773  ] =     26;
		rom[ 774  ] =   -188;
		rom[ 775  ] =    236;
		rom[ 776  ] =    -24;
		rom[ 777  ] =   -213;
		rom[ 778  ] =    190;
		rom[ 779  ] =     30;
		rom[ 780  ] =     88;
		rom[ 781  ] =    -73;
		rom[ 782  ] =   -152;
		rom[ 783  ] =     -1;
		rom[ 784  ] =    102;
		rom[ 785  ] =     38;
		rom[ 786  ] =    132;
		rom[ 787  ] =    -25;
		rom[ 788  ] =    210;
		rom[ 789  ] =   -108;
		rom[ 790  ] =    -63;
		rom[ 791  ] =     79;
		rom[ 792  ] =    137;
		rom[ 793  ] =    118;
		rom[ 794  ] =      0;
		rom[ 795  ] =   -201;
		rom[ 796  ] =    313;
		rom[ 797  ] =     97;
		rom[ 798  ] =     15;
		rom[ 799  ] =   -366;
		rom[ 800  ] =    -61;
		rom[ 801  ] =    -45;
		rom[ 802  ] =    387;
		rom[ 803  ] =   2254;
		rom[ 804  ] =    169;
		rom[ 805  ] =    101;
		rom[ 806  ] =    208;
		rom[ 807  ] =    -69;
		rom[ 808  ] =   -498;
		rom[ 809  ] =    -14;
		rom[ 810  ] =    474;
		rom[ 811  ] =    151;
		rom[ 812  ] =     47;
		rom[ 813  ] =    -82;
		rom[ 814  ] =   -117;
		rom[ 815  ] =    -23;
		rom[ 816  ] =   -227;
		rom[ 817  ] =    -60;
		rom[ 818  ] =    -29;
		rom[ 819  ] =   -184;
		rom[ 820  ] =    263;
		rom[ 821  ] =    -60;
		rom[ 822  ] =    184;
		rom[ 823  ] =     -4;
		rom[ 824  ] =    202;
		rom[ 825  ] =    119;
		rom[ 826  ] =    142;
		rom[ 827  ] =    -25;
		rom[ 828  ] =     63;
		rom[ 829  ] =     11;
		rom[ 830  ] =   -219;
		rom[ 831  ] =    -78;
		rom[ 832  ] =   -226;
		rom[ 833  ] =    230;
		rom[ 834  ] =    -97;
		rom[ 835  ] =      7;
		rom[ 836  ] =   -154;
		rom[ 837  ] =    -98;
		rom[ 838  ] =    112;
		rom[ 839  ] =    473;
		rom[ 840  ] =    -91;
		rom[ 841  ] =     54;
		rom[ 842  ] =    -15;
		rom[ 843  ] =    -10;
		rom[ 844  ] =     13;
		rom[ 845  ] =    154;
		rom[ 846  ] =    -56;
		rom[ 847  ] =    -11;
		rom[ 848  ] =   -157;
		rom[ 849  ] =   -142;
		rom[ 850  ] =     95;
		rom[ 851  ] =    143;
		rom[ 852  ] =    -54;
		rom[ 853  ] =     52;
		rom[ 854  ] =     14;
		rom[ 855  ] =    412;
		rom[ 856  ] =      0;
		rom[ 857  ] =     47;
		rom[ 858  ] =   -147;
		rom[ 859  ] =    -86;
		rom[ 860  ] =     60;
		rom[ 861  ] =    -21;
		rom[ 862  ] =     96;
		rom[ 863  ] =   -102;
		rom[ 864  ] =     -3;
		rom[ 865  ] =   -165;
		rom[ 866  ] =    115;
		rom[ 867  ] =    187;
		rom[ 868  ] =    162;
		rom[ 869  ] =    206;
		rom[ 870  ] =    -70;
		rom[ 871  ] =    328;
		rom[ 872  ] =    400;
		rom[ 873  ] =    -63;
		rom[ 874  ] =    -62;
		rom[ 875  ] =    -67;
		rom[ 876  ] =   -107;
		rom[ 877  ] =     36;
		rom[ 878  ] =   -110;
		rom[ 879  ] =     31;
		rom[ 880  ] =    -65;
		rom[ 881  ] =     85;
		rom[ 882  ] =    350;
		rom[ 883  ] =     97;
		rom[ 884  ] =   -160;
		rom[ 885  ] =   -319;
		rom[ 886  ] =    -69;
		rom[ 887  ] =    486;
		rom[ 888  ] =    639;
		rom[ 889  ] =   -188;
		rom[ 890  ] =    -42;
		rom[ 891  ] =    392;
		rom[ 892  ] =     56;
		rom[ 893  ] =      9;
		rom[ 894  ] =    136;
		rom[ 895  ] =   -136;
		rom[ 896  ] =     11;
		rom[ 897  ] =   -269;
		rom[ 898  ] =      8;
		rom[ 899  ] =     91;
		rom[ 900  ] =   -235;
		rom[ 901  ] =     27;
		rom[ 902  ] =     50;
		rom[ 903  ] =    -33;
		rom[ 904  ] =    150;
		rom[ 905  ] =  -1647;
		rom[ 906  ] =    -90;
		rom[ 907  ] =    -53;
		rom[ 908  ] =    -52;
		rom[ 909  ] =     88;
		rom[ 910  ] =     48;
		rom[ 911  ] =    -80;
		rom[ 912  ] =    263;
		rom[ 913  ] =    446;
		rom[ 914  ] =   -139;
		rom[ 915  ] =    -15;
		rom[ 916  ] =    -44;
		rom[ 917  ] =    -47;
		rom[ 918  ] =    106;
		rom[ 919  ] =     17;
		rom[ 920  ] =   -195;
		rom[ 921  ] =      1;
		rom[ 922  ] =    472;
		rom[ 923  ] =     65;
		rom[ 924  ] =    231;
		rom[ 925  ] =    -43;
		rom[ 926  ] =    508;
		rom[ 927  ] =    -22;
		rom[ 928  ] =     48;
		rom[ 929  ] =   -176;
		rom[ 930  ] =   -135;
		rom[ 931  ] =    -87;
		rom[ 932  ] =    -50;
		rom[ 933  ] =    -69;
		rom[ 934  ] =    -10;
		rom[ 935  ] =   -184;
		rom[ 936  ] =    159;
		rom[ 937  ] =     27;
		rom[ 938  ] =    -67;
		rom[ 939  ] =     25;
		rom[ 940  ] =    187;
		rom[ 941  ] =     16;
		rom[ 942  ] =      0;
		rom[ 943  ] =     29;
		rom[ 944  ] =   -204;
		rom[ 945  ] =   -102;
		rom[ 946  ] =    126;
		rom[ 947  ] =    189;
		rom[ 948  ] =    -13;
		rom[ 949  ] =    -99;
		rom[ 950  ] =     49;
		rom[ 951  ] =     53;
		rom[ 952  ] =    242;
		rom[ 953  ] =   -168;
		rom[ 954  ] =   -344;
		rom[ 955  ] =    182;
		rom[ 956  ] =    100;
		rom[ 957  ] =    -17;
		rom[ 958  ] =    100;
		rom[ 959  ] =   -348;
		rom[ 960  ] =     89;
		rom[ 961  ] =    -68;
		rom[ 962  ] =    133;
		rom[ 963  ] =     10;
		rom[ 964  ] =    226;
		rom[ 965  ] =   -435;
		rom[ 966  ] =    -32;
		rom[ 967  ] =    309;
		rom[ 968  ] =   -380;
		rom[ 969  ] =    202;
		rom[ 970  ] =    -48;
		rom[ 971  ] =    351;
		rom[ 972  ] =    331;
		rom[ 973  ] =   -138;
		rom[ 974  ] =     63;
		rom[ 975  ] =    224;
		rom[ 976  ] =     87;
		rom[ 977  ] =     32;
		rom[ 978  ] =   -153;
		rom[ 979  ] =    652;
		rom[ 980  ] =   -282;
		rom[ 981  ] =   -138;
		rom[ 982  ] =   -259;
		rom[ 983  ] =     30;
		rom[ 984  ] =    -39;
		rom[ 985  ] =   -535;
		rom[ 986  ] =    235;
		rom[ 987  ] =    -29;
		rom[ 988  ] =    127;
		rom[ 989  ] =    146;
		rom[ 990  ] =   -129;
		rom[ 991  ] =    -79;
		rom[ 992  ] =    -29;
		rom[ 993  ] =     33;
		rom[ 994  ] =   -178;
		rom[ 995  ] =    108;
		rom[ 996  ] =    131;
		rom[ 997  ] =   -295;
		rom[ 998  ] =    128;
		rom[ 999  ] =     -1;
		rom[ 1000 ] =     11;
		rom[ 1001 ] =    134;
		rom[ 1002 ] =    -59;
		rom[ 1003 ] =    155;
		rom[ 1004 ] =     11;
		rom[ 1005 ] =   -170;
		rom[ 1006 ] =   -101;
		rom[ 1007 ] =     41;
		rom[ 1008 ] =    -85;
		rom[ 1009 ] =     91;
		rom[ 1010 ] =   -152;
		rom[ 1011 ] =    -43;
		rom[ 1012 ] =    227;
		rom[ 1013 ] =     88;
		rom[ 1014 ] =      0;
		rom[ 1015 ] =     59;
		rom[ 1016 ] =    441;
		rom[ 1017 ] =    147;
		rom[ 1018 ] =    -16;
		rom[ 1019 ] =     85;
		rom[ 1020 ] =   -122;
		rom[ 1021 ] =    106;
		rom[ 1022 ] =     43;
		rom[ 1023 ] =     35;
		rom[ 1024 ] =     87;
		rom[ 1025 ] =    305;
		rom[ 1026 ] =     19;
		rom[ 1027 ] =      7;
		rom[ 1028 ] =      4;
		rom[ 1029 ] =    115;
		rom[ 1030 ] =   -133;
		rom[ 1031 ] =     92;
		rom[ 1032 ] =    -88;
		rom[ 1033 ] =     31;
		rom[ 1034 ] =     59;
		rom[ 1035 ] =    114;
		rom[ 1036 ] =     23;
		rom[ 1037 ] =    -40;
		rom[ 1038 ] =    -16;
		rom[ 1039 ] =    -92;
		rom[ 1040 ] =   -162;
		rom[ 1041 ] =    -71;
		rom[ 1042 ] =     36;
		rom[ 1043 ] =    -32;
		rom[ 1044 ] =    110;
		rom[ 1045 ] =    -84;
		rom[ 1046 ] =   -294;
		rom[ 1047 ] =   -110;
		rom[ 1048 ] =   -194;
		rom[ 1049 ] =   -446;
		rom[ 1050 ] =     55;
		rom[ 1051 ] =    -27;
		rom[ 1052 ] =    -16;
		rom[ 1053 ] =   -154;
		rom[ 1054 ] =     35;
		rom[ 1055 ] =   -131;
		rom[ 1056 ] =    239;
		rom[ 1057 ] =   -167;
		rom[ 1058 ] =    -81;
		rom[ 1059 ] =    -18;
		rom[ 1060 ] =     68;
		rom[ 1061 ] =     38;
		rom[ 1062 ] =    -80;
		rom[ 1063 ] =     44;
		rom[ 1064 ] =    155;
		rom[ 1065 ] =     67;
		rom[ 1066 ] =    -81;
		rom[ 1067 ] =     45;
		rom[ 1068 ] =     21;
		rom[ 1069 ] =    -45;
		rom[ 1070 ] =    -43;
		rom[ 1071 ] =    431;
		rom[ 1072 ] =    224;
		rom[ 1073 ] =     72;
		rom[ 1074 ] =   -127;
		rom[ 1075 ] =   -234;
		rom[ 1076 ] =    -46;
		rom[ 1077 ] =    125;
		rom[ 1078 ] =      7;
		rom[ 1079 ] =     46;
		rom[ 1080 ] =    333;
		rom[ 1081 ] =    219;
		rom[ 1082 ] =    -98;
		rom[ 1083 ] =     27;
		rom[ 1084 ] =   -132;
		rom[ 1085 ] =    155;
		rom[ 1086 ] =     63;
		rom[ 1087 ] =   -181;
		rom[ 1088 ] =    -94;
		rom[ 1089 ] =     79;
		rom[ 1090 ] =    425;
		rom[ 1091 ] =    -77;
		rom[ 1092 ] =    158;
		rom[ 1093 ] =     93;
		rom[ 1094 ] =   -128;
		rom[ 1095 ] =     39;
		rom[ 1096 ] =   -201;
		rom[ 1097 ] =   -161;
		rom[ 1098 ] =    196;
		rom[ 1099 ] =    210;
		rom[ 1100 ] =     58;
		rom[ 1101 ] =   -375;
		rom[ 1102 ] =     26;
		rom[ 1103 ] =    146;
		rom[ 1104 ] =    207;
		rom[ 1105 ] =    -59;
		rom[ 1106 ] =   -158;
		rom[ 1107 ] =   -165;
		rom[ 1108 ] =     97;
		rom[ 1109 ] =     35;
		rom[ 1110 ] =   -544;
		rom[ 1111 ] =     40;
		rom[ 1112 ] =     20;
		rom[ 1113 ] =   -250;
		rom[ 1114 ] =     -1;
		rom[ 1115 ] =     13;
		rom[ 1116 ] =     86;
		rom[ 1117 ] =     30;
		rom[ 1118 ] =    101;
		rom[ 1119 ] =   -145;
		rom[ 1120 ] =     81;
		rom[ 1121 ] =     61;
		rom[ 1122 ] =    -94;
		rom[ 1123 ] =    -76;
		rom[ 1124 ] =   1846;
		rom[ 1125 ] =     48;
		rom[ 1126 ] =   -101;
		rom[ 1127 ] =   -183;
		rom[ 1128 ] =    -59;
		rom[ 1129 ] =   -100;
		rom[ 1130 ] =     94;
		rom[ 1131 ] =   -102;
		rom[ 1132 ] =      4;
		rom[ 1133 ] =     63;
		rom[ 1134 ] =   -109;
		rom[ 1135 ] =      5;
		rom[ 1136 ] =     -2;
		rom[ 1137 ] =   -130;
		rom[ 1138 ] =    -20;
		rom[ 1139 ] =    127;
		rom[ 1140 ] =   -137;
		rom[ 1141 ] =     49;
		rom[ 1142 ] =   -142;
		rom[ 1143 ] =     40;
		rom[ 1144 ] =    244;
		rom[ 1145 ] =   -267;
		rom[ 1146 ] =   -380;
		rom[ 1147 ] =   -168;
		rom[ 1148 ] =     87;
		rom[ 1149 ] =   -104;
		rom[ 1150 ] =   -168;
		rom[ 1151 ] =    -72;
		rom[ 1152 ] =     36;
		rom[ 1153 ] =    -47;
		rom[ 1154 ] =    -30;
		rom[ 1155 ] =      3;
		rom[ 1156 ] =   -125;
		rom[ 1157 ] =    -77;
		rom[ 1158 ] =    -33;
		rom[ 1159 ] =   -142;
		rom[ 1160 ] =     77;
		rom[ 1161 ] =    -77;
		rom[ 1162 ] =   -364;
		rom[ 1163 ] =     28;
		rom[ 1164 ] =   -115;
		rom[ 1165 ] =     -1;
		rom[ 1166 ] =   -443;
		rom[ 1167 ] =     65;
		rom[ 1168 ] =     35;
		rom[ 1169 ] =   -103;
		rom[ 1170 ] =    -55;
		rom[ 1171 ] =    -31;
		rom[ 1172 ] =    293;
		rom[ 1173 ] =    -55;
		rom[ 1174 ] =     12;
		rom[ 1175 ] =   -208;
		rom[ 1176 ] =    -36;
		rom[ 1177 ] =    877;
		rom[ 1178 ] =     57;
		rom[ 1179 ] =    174;
		rom[ 1180 ] =     81;
		rom[ 1181 ] =   -137;
		rom[ 1182 ] =    260;
		rom[ 1183 ] =     89;
		rom[ 1184 ] =   -321;
		rom[ 1185 ] =     58;
		rom[ 1186 ] =   -275;
		rom[ 1187 ] =    534;
		rom[ 1188 ] =   -189;
		rom[ 1189 ] =   -122;
		rom[ 1190 ] =     -1;
		rom[ 1191 ] =    -91;
		rom[ 1192 ] =     -6;
		rom[ 1193 ] =     49;
		rom[ 1194 ] =     99;
		rom[ 1195 ] =   -193;
		rom[ 1196 ] =   -101;
		rom[ 1197 ] =     89;
		rom[ 1198 ] =    770;
		rom[ 1199 ] =   -318;
		rom[ 1200 ] =   -199;
		rom[ 1201 ] =    -70;
		rom[ 1202 ] =    -11;
		rom[ 1203 ] =   -404;
		rom[ 1204 ] =    -89;
		rom[ 1205 ] =    250;
		rom[ 1206 ] =   -100;
		rom[ 1207 ] =    138;
		rom[ 1208 ] =    156;
		rom[ 1209 ] =    -82;
		rom[ 1210 ] =    101;
		rom[ 1211 ] =    -99;
		rom[ 1212 ] =   -108;
		rom[ 1213 ] =    -14;
		rom[ 1214 ] =    438;
		rom[ 1215 ] =    184;
		rom[ 1216 ] =    181;
		rom[ 1217 ] =      4;
		rom[ 1218 ] =    292;
		rom[ 1219 ] =    146;
		rom[ 1220 ] =    -85;
		rom[ 1221 ] =   1741;
		rom[ 1222 ] =     46;
		rom[ 1223 ] =    -62;
		rom[ 1224 ] =    -62;
		rom[ 1225 ] =    -77;
		rom[ 1226 ] =    -13;
		rom[ 1227 ] =    381;
		rom[ 1228 ] =    -51;
		rom[ 1229 ] =   -110;
		rom[ 1230 ] =    -96;
		rom[ 1231 ] =    -58;
		rom[ 1232 ] =    115;
		rom[ 1233 ] =    208;
		rom[ 1234 ] =     47;
		rom[ 1235 ] =    -60;
		rom[ 1236 ] =    935;
		rom[ 1237 ] =    454;
		rom[ 1238 ] =     13;
		rom[ 1239 ] =    349;
		rom[ 1240 ] =     90;
		rom[ 1241 ] =    -64;
		rom[ 1242 ] =   1356;
		rom[ 1243 ] =     36;
		rom[ 1244 ] =    188;
		rom[ 1245 ] =   -154;
		rom[ 1246 ] =   -335;
		rom[ 1247 ] =    891;
		rom[ 1248 ] =     60;
		rom[ 1249 ] =    214;
		rom[ 1250 ] =     37;
		rom[ 1251 ] =     32;
		rom[ 1252 ] =   -106;
		rom[ 1253 ] =    -12;
		rom[ 1254 ] =    234;
		rom[ 1255 ] =    -25;
		rom[ 1256 ] =   -165;
		rom[ 1257 ] =    -83;
		rom[ 1258 ] =    -70;
		rom[ 1259 ] =    -99;
		rom[ 1260 ] =    232;
		rom[ 1261 ] =      1;
		rom[ 1262 ] =     40;
		rom[ 1263 ] =   -215;
		rom[ 1264 ] =    -56;
		rom[ 1265 ] =   -124;
		rom[ 1266 ] =  -1230;
		rom[ 1267 ] =   -147;
		rom[ 1268 ] =   -225;
		rom[ 1269 ] =    138;
		rom[ 1270 ] =    -33;
		rom[ 1271 ] =    -22;
		rom[ 1272 ] =     12;
		rom[ 1273 ] =    219;
		rom[ 1274 ] =   -513;
		rom[ 1275 ] =    379;
		rom[ 1276 ] =    157;
		rom[ 1277 ] =     -8;
		rom[ 1278 ] =     39;
		rom[ 1279 ] =     98;
		rom[ 1280 ] =    -73;
		rom[ 1281 ] =    -43;
		rom[ 1282 ] =    -29;
		rom[ 1283 ] =     98;
		rom[ 1284 ] =    -75;
		rom[ 1285 ] =     64;
		rom[ 1286 ] =   -199;
		rom[ 1287 ] =     27;
		rom[ 1288 ] =     40;
		rom[ 1289 ] =     60;
		rom[ 1290 ] =    397;
		rom[ 1291 ] =    197;
		rom[ 1292 ] =     40;
		rom[ 1293 ] =   -163;
		rom[ 1294 ] =     93;
		rom[ 1295 ] =     27;
		rom[ 1296 ] =    244;
		rom[ 1297 ] =     28;
		rom[ 1298 ] =     64;
		rom[ 1299 ] =   -203;
		rom[ 1300 ] =    214;
		rom[ 1301 ] =     91;
		rom[ 1302 ] =    168;
		rom[ 1303 ] =    -88;
		rom[ 1304 ] =   -339;
		rom[ 1305 ] =     34;
		rom[ 1306 ] =    323;
		rom[ 1307 ] =   -369;
		rom[ 1308 ] =   -119;
		rom[ 1309 ] =     28;
		rom[ 1310 ] =    -33;
		rom[ 1311 ] =     80;
		rom[ 1312 ] =    -60;
		rom[ 1313 ] =    103;
		rom[ 1314 ] =    -64;
		rom[ 1315 ] =    120;
		rom[ 1316 ] =    -34;
		rom[ 1317 ] =    100;
		rom[ 1318 ] =   -138;
		rom[ 1319 ] =     -8;
		rom[ 1320 ] =    124;
		rom[ 1321 ] =     16;
		rom[ 1322 ] =    113;
		rom[ 1323 ] =     32;
		rom[ 1324 ] =    180;
		rom[ 1325 ] =   -132;
		rom[ 1326 ] =     85;
		rom[ 1327 ] =    103;
		rom[ 1328 ] =     26;
		rom[ 1329 ] =   -239;
		rom[ 1330 ] =    130;
		rom[ 1331 ] =   -124;
		rom[ 1332 ] =     61;
		rom[ 1333 ] =   -200;
		rom[ 1334 ] =    340;
		rom[ 1335 ] =     97;
		rom[ 1336 ] =     67;
		rom[ 1337 ] =    -48;
		rom[ 1338 ] =      0;
		rom[ 1339 ] =     78;
		rom[ 1340 ] =    -41;
		rom[ 1341 ] =    -57;
		rom[ 1342 ] =   -422;
		rom[ 1343 ] =   -391;
		rom[ 1344 ] =   -169;
		rom[ 1345 ] =      9;
		rom[ 1346 ] =    439;
		rom[ 1347 ] =     13;
		rom[ 1348 ] =    119;
		rom[ 1349 ] =     46;
		rom[ 1350 ] =    -49;
		rom[ 1351 ] =    -52;
		rom[ 1352 ] =    100;
		rom[ 1353 ] =    188;
		rom[ 1354 ] =   -111;
		rom[ 1355 ] =    164;
		rom[ 1356 ] =     94;
		rom[ 1357 ] =    -97;
		rom[ 1358 ] =    317;
		rom[ 1359 ] =    -54;
		rom[ 1360 ] =    -88;
		rom[ 1361 ] =   -292;
		rom[ 1362 ] =    -22;
		rom[ 1363 ] =    109;
		rom[ 1364 ] =   -161;
		rom[ 1365 ] =    106;
		rom[ 1366 ] =    200;
		rom[ 1367 ] =    151;
		rom[ 1368 ] =    323;
		rom[ 1369 ] =    118;
		rom[ 1370 ] =     25;
		rom[ 1371 ] =   -269;
		rom[ 1372 ] =   -282;
		rom[ 1373 ] =   -477;
		rom[ 1374 ] =     -5;
		rom[ 1375 ] =   -182;
		rom[ 1376 ] =    209;
		rom[ 1377 ] =   -129;
		rom[ 1378 ] =     86;
		rom[ 1379 ] =   -566;
		rom[ 1380 ] =    213;
		rom[ 1381 ] =    106;
		rom[ 1382 ] =    -49;
		rom[ 1383 ] =    -99;
		rom[ 1384 ] =   -103;
		rom[ 1385 ] =     51;
		rom[ 1386 ] =    234;
		rom[ 1387 ] =     68;
		rom[ 1388 ] =    -93;
		rom[ 1389 ] =      0;
		rom[ 1390 ] =    -31;
		rom[ 1391 ] =    385;
		rom[ 1392 ] =   -255;
		rom[ 1393 ] =     71;
		rom[ 1394 ] =    -90;
		rom[ 1395 ] =    -42;
		rom[ 1396 ] =    -38;
		rom[ 1397 ] =   -118;
		rom[ 1398 ] =    -86;
		rom[ 1399 ] =   -151;
		rom[ 1400 ] =     43;
		rom[ 1401 ] =    670;
		rom[ 1402 ] =    388;
		rom[ 1403 ] =    144;
		rom[ 1404 ] =     52;
		rom[ 1405 ] =    569;
		rom[ 1406 ] =     48;
		rom[ 1407 ] =    -40;
		rom[ 1408 ] =    -24;
		rom[ 1409 ] =     -5;
		rom[ 1410 ] =    132;
		rom[ 1411 ] =    -57;
		rom[ 1412 ] =      4;
		rom[ 1413 ] =      0;
		rom[ 1414 ] =     -1;
		rom[ 1415 ] =     16;
		rom[ 1416 ] =     58;
		rom[ 1417 ] =   -226;
		rom[ 1418 ] =    383;
		rom[ 1419 ] =    109;
		rom[ 1420 ] =     15;
		rom[ 1421 ] =   -130;
		rom[ 1422 ] =    -92;
		rom[ 1423 ] =    103;
		rom[ 1424 ] =   -127;
		rom[ 1425 ] =   -108;
		rom[ 1426 ] =    -56;
		rom[ 1427 ] =   -257;
		rom[ 1428 ] =   -183;
		rom[ 1429 ] =    -83;
		rom[ 1430 ] =    -32;
		rom[ 1431 ] =     35;
		rom[ 1432 ] =   -111;
		rom[ 1433 ] =    -67;
		rom[ 1434 ] =    -56;
		rom[ 1435 ] =    119;
		rom[ 1436 ] =    153;
		rom[ 1437 ] =   -102;
		rom[ 1438 ] =   -261;
		rom[ 1439 ] =    -38;
		rom[ 1440 ] =     -3;
		rom[ 1441 ] =    -89;
		rom[ 1442 ] =    -73;
		rom[ 1443 ] =   -101;
		rom[ 1444 ] =    643;
		rom[ 1445 ] =    282;
		rom[ 1446 ] =    -45;
		rom[ 1447 ] =    -56;
		rom[ 1448 ] =   -126;
		rom[ 1449 ] =     87;
		rom[ 1450 ] =    381;
		rom[ 1451 ] =    121;
		rom[ 1452 ] =      0;
		rom[ 1453 ] =   -172;
		rom[ 1454 ] =    -92;
		rom[ 1455 ] =    -52;
		rom[ 1456 ] =    114;
		rom[ 1457 ] =   -113;
		rom[ 1458 ] =    -25;
		rom[ 1459 ] =    -83;
		rom[ 1460 ] =    -50;
		rom[ 1461 ] =   -165;
		rom[ 1462 ] =    121;
		rom[ 1463 ] =     28;
		rom[ 1464 ] =     66;
		rom[ 1465 ] =    205;
		rom[ 1466 ] =      8;
		rom[ 1467 ] =    102;
		rom[ 1468 ] =    -64;
		rom[ 1469 ] =    152;
		rom[ 1470 ] =   -324;
		rom[ 1471 ] =    -70;
		rom[ 1472 ] =    134;
		rom[ 1473 ] =   -481;
		rom[ 1474 ] =    493;
		rom[ 1475 ] =     17;
		rom[ 1476 ] =   -297;
		rom[ 1477 ] =    725;
		rom[ 1478 ] =     34;
		rom[ 1479 ] =    -53;
		rom[ 1480 ] =     77;
		rom[ 1481 ] =     87;
		rom[ 1482 ] =    259;
		rom[ 1483 ] =   -132;
		rom[ 1484 ] =    -96;
		rom[ 1485 ] =     76;
		rom[ 1486 ] =    127;
		rom[ 1487 ] =    -45;
		rom[ 1488 ] =    -52;
		rom[ 1489 ] =    -52;
		rom[ 1490 ] =    281;
		rom[ 1491 ] =     21;
		rom[ 1492 ] =   -158;
		rom[ 1493 ] =     25;
		rom[ 1494 ] =    717;
		rom[ 1495 ] =    476;
		rom[ 1496 ] =    -94;
		rom[ 1497 ] =   -210;
		rom[ 1498 ] =    920;
		rom[ 1499 ] =     38;
		rom[ 1500 ] =   -485;
		rom[ 1501 ] =    154;
		rom[ 1502 ] =     90;
		rom[ 1503 ] =   -148;
		rom[ 1504 ] =   -540;
		rom[ 1505 ] =   -170;
		rom[ 1506 ] =   -135;
		rom[ 1507 ] =     64;
		rom[ 1508 ] =   -161;
		rom[ 1509 ] =   -277;
		rom[ 1510 ] =   -109;
		rom[ 1511 ] =    163;
		rom[ 1512 ] =    412;
		rom[ 1513 ] =   -331;
		rom[ 1514 ] =    -87;
		rom[ 1515 ] =    -43;
		rom[ 1516 ] =      3;
		rom[ 1517 ] =     14;
		rom[ 1518 ] =     77;
		rom[ 1519 ] =   -104;
		rom[ 1520 ] =    -16;
		rom[ 1521 ] =     -3;
		rom[ 1522 ] =   -202;
		rom[ 1523 ] =     47;
		rom[ 1524 ] =    141;
		rom[ 1525 ] =    -33;
		rom[ 1526 ] =    -91;
		rom[ 1527 ] =   -126;
		rom[ 1528 ] =    179;
		rom[ 1529 ] =    176;
		rom[ 1530 ] =    111;
		rom[ 1531 ] =     38;
		rom[ 1532 ] =    386;
		rom[ 1533 ] =    697;
		rom[ 1534 ] =   -193;
		rom[ 1535 ] =    458;
		rom[ 1536 ] =    -58;
		rom[ 1537 ] =    139;
		rom[ 1538 ] =     88;
		rom[ 1539 ] =     89;
		rom[ 1540 ] =    337;
		rom[ 1541 ] =    346;
		rom[ 1542 ] =   -225;
		rom[ 1543 ] =   -265;
		rom[ 1544 ] =    -93;
		rom[ 1545 ] =    224;
		rom[ 1546 ] =      0;
		rom[ 1547 ] =    402;
		rom[ 1548 ] =    -29;
		rom[ 1549 ] =    205;
		rom[ 1550 ] =    -23;
		rom[ 1551 ] =     57;
		rom[ 1552 ] =     87;
		rom[ 1553 ] =   -119;
		rom[ 1554 ] =      1;
		rom[ 1555 ] =      7;
		rom[ 1556 ] =     35;
		rom[ 1557 ] =    260;
		rom[ 1558 ] =   -114;
		rom[ 1559 ] =    200;
		rom[ 1560 ] =   -120;
		rom[ 1561 ] =    508;
		rom[ 1562 ] =     32;
		rom[ 1563 ] =    124;
		rom[ 1564 ] =    103;
		rom[ 1565 ] =     41;
		rom[ 1566 ] =    -68;
		rom[ 1567 ] =    -11;
		rom[ 1568 ] =    173;
		rom[ 1569 ] =   -198;
		rom[ 1570 ] =    118;
		rom[ 1571 ] =   -164;
		rom[ 1572 ] =   -168;
		rom[ 1573 ] =     48;
		rom[ 1574 ] =    -87;
		rom[ 1575 ] =    -97;
		rom[ 1576 ] =     73;
		rom[ 1577 ] =   -178;
		rom[ 1578 ] =    -37;
		rom[ 1579 ] =    194;
		rom[ 1580 ] =    -58;
		rom[ 1581 ] =     15;
		rom[ 1582 ] =     14;
		rom[ 1583 ] =   -119;
		rom[ 1584 ] =    -26;
		rom[ 1585 ] =   -123;
		rom[ 1586 ] =     32;
		rom[ 1587 ] =     36;
		rom[ 1588 ] =    393;
		rom[ 1589 ] =   -134;
		rom[ 1590 ] =    -54;
		rom[ 1591 ] =     62;
		rom[ 1592 ] =     49;
		rom[ 1593 ] =   -312;
		rom[ 1594 ] =    -49;
		rom[ 1595 ] =     89;
		rom[ 1596 ] =    -11;
		rom[ 1597 ] =   -199;
		rom[ 1598 ] =    -42;
		rom[ 1599 ] =    -27;
		rom[ 1600 ] =     35;
		rom[ 1601 ] =     81;
		rom[ 1602 ] =     90;
		rom[ 1603 ] =   -213;
		rom[ 1604 ] =     80;
		rom[ 1605 ] =     94;
		rom[ 1606 ] =    -61;
		rom[ 1607 ] =   -204;
		rom[ 1608 ] =   -283;
		rom[ 1609 ] =     19;
		rom[ 1610 ] =   -138;
		rom[ 1611 ] =    -66;
		rom[ 1612 ] =   -205;
		rom[ 1613 ] =    233;
		rom[ 1614 ] =    167;
		rom[ 1615 ] =    -12;
		rom[ 1616 ] =   -133;
		rom[ 1617 ] =    403;
		rom[ 1618 ] =   -156;
		rom[ 1619 ] =   -188;
		rom[ 1620 ] =   -489;
		rom[ 1621 ] =   -493;
		rom[ 1622 ] =    289;
		rom[ 1623 ] =     34;
		rom[ 1624 ] =     93;
		rom[ 1625 ] =      2;
		rom[ 1626 ] =    141;
		rom[ 1627 ] =    -18;
		rom[ 1628 ] =     96;
		rom[ 1629 ] =     52;
		rom[ 1630 ] =    -46;
		rom[ 1631 ] =   -170;
		rom[ 1632 ] =   -382;
		rom[ 1633 ] =   -111;
		rom[ 1634 ] =    -89;
		rom[ 1635 ] =    -39;
		rom[ 1636 ] =    284;
		rom[ 1637 ] =    127;
		rom[ 1638 ] =   -203;
		rom[ 1639 ] =    -83;
		rom[ 1640 ] =    -62;
		rom[ 1641 ] =   -207;
		rom[ 1642 ] =    -84;
		rom[ 1643 ] =   -126;
		rom[ 1644 ] =    -18;
		rom[ 1645 ] =   -187;
		rom[ 1646 ] =     68;
		rom[ 1647 ] =     13;
		rom[ 1648 ] =    100;
		rom[ 1649 ] =   -326;
		rom[ 1650 ] =    182;
		rom[ 1651 ] =   -513;
		rom[ 1652 ] =     73;
		rom[ 1653 ] =     78;
		rom[ 1654 ] =    163;
		rom[ 1655 ] =     55;
		rom[ 1656 ] =     66;
		rom[ 1657 ] =     45;
		rom[ 1658 ] =    160;
		rom[ 1659 ] =    -39;
		rom[ 1660 ] =    114;
		rom[ 1661 ] =    -96;
		rom[ 1662 ] =    110;
		rom[ 1663 ] =      1;
		rom[ 1664 ] =   -168;
		rom[ 1665 ] =     27;
		rom[ 1666 ] =    196;
		rom[ 1667 ] =    -12;
		rom[ 1668 ] =    -35;
		rom[ 1669 ] =    -30;
		rom[ 1670 ] =     -7;
		rom[ 1671 ] =   -353;
		rom[ 1672 ] =    191;
		rom[ 1673 ] =      0;
		rom[ 1674 ] =    -66;
		rom[ 1675 ] =    187;
		rom[ 1676 ] =   -112;
		rom[ 1677 ] =   -113;
		rom[ 1678 ] =     31;
		rom[ 1679 ] =     -2;
		rom[ 1680 ] =    452;
		rom[ 1681 ] =    281;
		rom[ 1682 ] =      7;
		rom[ 1683 ] =    787;
		rom[ 1684 ] =    644;
		rom[ 1685 ] =   -202;
		rom[ 1686 ] =    212;
		rom[ 1687 ] =    204;
		rom[ 1688 ] =   -174;
		rom[ 1689 ] =   -153;
		rom[ 1690 ] =   -152;
		rom[ 1691 ] =     57;
		rom[ 1692 ] =     -1;
		rom[ 1693 ] =    131;
		rom[ 1694 ] =    -17;
		rom[ 1695 ] =     40;
		rom[ 1696 ] =    382;
		rom[ 1697 ] =     70;
		rom[ 1698 ] =     34;
		rom[ 1699 ] =    -57;
		rom[ 1700 ] =    -31;
		rom[ 1701 ] =    114;
		rom[ 1702 ] =    -77;
		rom[ 1703 ] =    -76;
		rom[ 1704 ] =   -149;
		rom[ 1705 ] =    132;
		rom[ 1706 ] =    244;
		rom[ 1707 ] =     40;
		rom[ 1708 ] =   -144;
		rom[ 1709 ] =     11;
		rom[ 1710 ] =     33;
		rom[ 1711 ] =    364;
		rom[ 1712 ] =   -123;
		rom[ 1713 ] =    -89;
		rom[ 1714 ] =    154;
		rom[ 1715 ] =     11;
		rom[ 1716 ] =    -43;
		rom[ 1717 ] =    531;
		rom[ 1718 ] =    -72;
		rom[ 1719 ] =   -315;
		rom[ 1720 ] =    -78;
		rom[ 1721 ] =   -209;
		rom[ 1722 ] =      8;
		rom[ 1723 ] =    104;
		rom[ 1724 ] =    -97;
		rom[ 1725 ] =    -26;
		rom[ 1726 ] =   -154;
		rom[ 1727 ] =    886;
		rom[ 1728 ] =    -54;
		rom[ 1729 ] =    291;
		rom[ 1730 ] =    229;
		rom[ 1731 ] =    165;
		rom[ 1732 ] =    258;
		rom[ 1733 ] =     42;
		rom[ 1734 ] =    256;
		rom[ 1735 ] =   -161;
		rom[ 1736 ] =    -22;
		rom[ 1737 ] =    441;
		rom[ 1738 ] =     69;
		rom[ 1739 ] =    127;
		rom[ 1740 ] =    -94;
		rom[ 1741 ] =    -45;
		rom[ 1742 ] =    -19;
		rom[ 1743 ] =    -71;
		rom[ 1744 ] =     77;
		rom[ 1745 ] =     29;
		rom[ 1746 ] =     77;
		rom[ 1747 ] =    127;
		rom[ 1748 ] =     85;
		rom[ 1749 ] =     46;
		rom[ 1750 ] =   -233;
		rom[ 1751 ] =    295;
		rom[ 1752 ] =    -81;
		rom[ 1753 ] =    -68;
		rom[ 1754 ] =   -163;
		rom[ 1755 ] =    110;
		rom[ 1756 ] =    -16;
		rom[ 1757 ] =     93;
		rom[ 1758 ] =   -282;
		rom[ 1759 ] =    176;
		rom[ 1760 ] =     35;
		rom[ 1761 ] =     59;
		rom[ 1762 ] =    -47;
		rom[ 1763 ] =   -449;
		rom[ 1764 ] =    185;
		rom[ 1765 ] =   -110;
		rom[ 1766 ] =     73;
		rom[ 1767 ] =    206;
		rom[ 1768 ] =   -122;
		rom[ 1769 ] =    155;
		rom[ 1770 ] =    760;
		rom[ 1771 ] =    -16;
		rom[ 1772 ] =     41;
		rom[ 1773 ] =    -47;
		rom[ 1774 ] =    -26;
		rom[ 1775 ] =     43;
		rom[ 1776 ] =    -83;
		rom[ 1777 ] =      9;
		rom[ 1778 ] =     -6;
		rom[ 1779 ] =     35;
		rom[ 1780 ] =    -99;
		rom[ 1781 ] =    304;
		rom[ 1782 ] =     69;
		rom[ 1783 ] =   -100;
		rom[ 1784 ] =    123;
		rom[ 1785 ] =     49;
		rom[ 1786 ] =    355;
		rom[ 1787 ] =   -173;
		rom[ 1788 ] =    -10;
		rom[ 1789 ] =   -232;
		rom[ 1790 ] =     96;
		rom[ 1791 ] =    -85;
		rom[ 1792 ] =     29;
		rom[ 1793 ] =   1399;
		rom[ 1794 ] =     25;
		rom[ 1795 ] =    133;
		rom[ 1796 ] =      0;
		rom[ 1797 ] =      2;
		rom[ 1798 ] =    223;
		rom[ 1799 ] =    -41;
		rom[ 1800 ] =    -77;
		rom[ 1801 ] =    -21;
		rom[ 1802 ] =    -44;
		rom[ 1803 ] =   -204;
		rom[ 1804 ] =     49;
		rom[ 1805 ] =     -9;
		rom[ 1806 ] =     12;
		rom[ 1807 ] =     16;
		rom[ 1808 ] =    -30;
		rom[ 1809 ] =    212;
		rom[ 1810 ] =     75;
		rom[ 1811 ] =    716;
		rom[ 1812 ] =    221;
		rom[ 1813 ] =  -1312;
		rom[ 1814 ] =   -110;
		rom[ 1815 ] =    317;
		rom[ 1816 ] =     97;
		rom[ 1817 ] =     47;
		rom[ 1818 ] =    133;
		rom[ 1819 ] =   -181;
		rom[ 1820 ] =   -239;
		rom[ 1821 ] =     79;
		rom[ 1822 ] =   -183;
		rom[ 1823 ] =   -247;
		rom[ 1824 ] =     47;
		rom[ 1825 ] =    114;
		rom[ 1826 ] =    267;
		rom[ 1827 ] =     39;
		rom[ 1828 ] =     10;
		rom[ 1829 ] =    130;
		rom[ 1830 ] =    135;
		rom[ 1831 ] =    194;
		rom[ 1832 ] =    -80;
		rom[ 1833 ] =   -224;
		rom[ 1834 ] =    -92;
		rom[ 1835 ] =    438;
		rom[ 1836 ] =   -149;
		rom[ 1837 ] =     57;
		rom[ 1838 ] =     85;
		rom[ 1839 ] =    201;
		rom[ 1840 ] =    148;
		rom[ 1841 ] =    168;
		rom[ 1842 ] =     64;
		rom[ 1843 ] =    -66;
		rom[ 1844 ] =    -12;
		rom[ 1845 ] =   -564;
		rom[ 1846 ] =    -39;
		rom[ 1847 ] =   -101;
		rom[ 1848 ] =   -571;
		rom[ 1849 ] =   -336;
		rom[ 1850 ] =     15;
		rom[ 1851 ] =    -27;
		rom[ 1852 ] =    -65;
		rom[ 1853 ] =   -208;
		rom[ 1854 ] =     68;
		rom[ 1855 ] =     65;
		rom[ 1856 ] =     14;
		rom[ 1857 ] =   -352;
		rom[ 1858 ] =    135;
		rom[ 1859 ] =    -16;
		rom[ 1860 ] =    -98;
		rom[ 1861 ] =     35;
		rom[ 1862 ] =   -113;
		rom[ 1863 ] =   -796;
		rom[ 1864 ] =   -445;
		rom[ 1865 ] =    -79;
		rom[ 1866 ] =     12;
		rom[ 1867 ] =    242;
		rom[ 1868 ] =   -222;
		rom[ 1869 ] =   -161;
		rom[ 1870 ] =    337;
		rom[ 1871 ] =    -30;
		rom[ 1872 ] =     30;
		rom[ 1873 ] =     28;
		rom[ 1874 ] =    -63;
		rom[ 1875 ] =    -11;
		rom[ 1876 ] =   -289;
		rom[ 1877 ] =    -47;
		rom[ 1878 ] =      2;
		rom[ 1879 ] =   -151;
		rom[ 1880 ] =   -133;
		rom[ 1881 ] =   -306;
		rom[ 1882 ] =    169;
		rom[ 1883 ] =   -118;
		rom[ 1884 ] =    189;
		rom[ 1885 ] =   1041;
		rom[ 1886 ] =      9;
		rom[ 1887 ] =   -339;
		rom[ 1888 ] =    -46;
		rom[ 1889 ] =   -528;
		rom[ 1890 ] =    157;
		rom[ 1891 ] =    417;
		rom[ 1892 ] =    -78;
		rom[ 1893 ] =   -248;
		rom[ 1894 ] =    101;
		rom[ 1895 ] =    109;
		rom[ 1896 ] =     61;
		rom[ 1897 ] =    107;
		rom[ 1898 ] =   -153;
		rom[ 1899 ] =    -21;
		rom[ 1900 ] =     72;
		rom[ 1901 ] =   -139;
		rom[ 1902 ] =    -65;
		rom[ 1903 ] =     80;
		rom[ 1904 ] =   -424;
		rom[ 1905 ] =    -78;
		rom[ 1906 ] =    -52;
		rom[ 1907 ] =    -66;
		rom[ 1908 ] =   -522;
		rom[ 1909 ] =     78;
		rom[ 1910 ] =    133;
		rom[ 1911 ] =     38;
		rom[ 1912 ] =     20;
		rom[ 1913 ] =    169;
		rom[ 1914 ] =   -312;
		rom[ 1915 ] =   -298;
		rom[ 1916 ] =    244;
		rom[ 1917 ] =     83;
		rom[ 1918 ] =   -328;
		rom[ 1919 ] =    -73;
		rom[ 1920 ] =     46;
		rom[ 1921 ] =   -104;
		rom[ 1922 ] =     -3;
		rom[ 1923 ] =    -59;
		rom[ 1924 ] =     35;
		rom[ 1925 ] =    224;
		rom[ 1926 ] =   -443;
		rom[ 1927 ] =     94;
		rom[ 1928 ] =     11;
		rom[ 1929 ] =     -8;
		rom[ 1930 ] =    -92;
		rom[ 1931 ] =    340;
		rom[ 1932 ] =    -27;
		rom[ 1933 ] =    313;
		rom[ 1934 ] =     22;
		rom[ 1935 ] =    -42;
		rom[ 1936 ] =    113;
		rom[ 1937 ] =    -95;
		rom[ 1938 ] =   -227;
		rom[ 1939 ] =   -166;
		rom[ 1940 ] =    -30;
		rom[ 1941 ] =     69;
		rom[ 1942 ] =   -151;
		rom[ 1943 ] =    -80;
		rom[ 1944 ] =    -96;
		rom[ 1945 ] =   -177;
		rom[ 1946 ] =    -90;
		rom[ 1947 ] =     67;
		rom[ 1948 ] =   -134;
		rom[ 1949 ] =    292;
		rom[ 1950 ] =      3;
		rom[ 1951 ] =    -34;
		rom[ 1952 ] =    -70;
		rom[ 1953 ] =    -76;
		rom[ 1954 ] =    -37;
		rom[ 1955 ] =     75;
		rom[ 1956 ] =   -206;
		rom[ 1957 ] =    -96;
		rom[ 1958 ] =   -111;
		rom[ 1959 ] =     26;
		rom[ 1960 ] =     95;
		rom[ 1961 ] =     53;
		rom[ 1962 ] =    -27;
		rom[ 1963 ] =    -92;
		rom[ 1964 ] =   -261;
		rom[ 1965 ] =   -204;
		rom[ 1966 ] =     27;
		rom[ 1967 ] =   -228;
		rom[ 1968 ] =   1308;
		rom[ 1969 ] =    331;
		rom[ 1970 ] =    -61;
		rom[ 1971 ] =    191;
		rom[ 1972 ] =     24;
		rom[ 1973 ] =   -140;
		rom[ 1974 ] =   -143;
		rom[ 1975 ] =     12;
		rom[ 1976 ] =    -57;
		rom[ 1977 ] =    -27;
		rom[ 1978 ] =   -216;
		rom[ 1979 ] =     -8;
		rom[ 1980 ] =     75;
		rom[ 1981 ] =     51;
		rom[ 1982 ] =     52;
		rom[ 1983 ] =    -73;
		rom[ 1984 ] =      7;
		rom[ 1985 ] =    -60;
		rom[ 1986 ] =    -61;
		rom[ 1987 ] =     59;
		rom[ 1988 ] =    -44;
		rom[ 1989 ] =    -37;
		rom[ 1990 ] =     18;
		rom[ 1991 ] =     96;
		rom[ 1992 ] =    130;
		rom[ 1993 ] =    -75;
		rom[ 1994 ] =     80;
		rom[ 1995 ] =   1685;
		rom[ 1996 ] =   -170;
		rom[ 1997 ] =    -42;
		rom[ 1998 ] =     50;
		rom[ 1999 ] =    -35;
		rom[ 2000 ] =     66;
		rom[ 2001 ] =    -42;
		rom[ 2002 ] =    -50;
		rom[ 2003 ] =   -206;
		rom[ 2004 ] =    202;
		rom[ 2005 ] =   -168;
		rom[ 2006 ] =      4;
		rom[ 2007 ] =   -205;
		rom[ 2008 ] =    -35;
		rom[ 2009 ] =   -205;
		rom[ 2010 ] =    418;
		rom[ 2011 ] =    -58;
		rom[ 2012 ] =     42;
		rom[ 2013 ] =    -48;
		rom[ 2014 ] =    295;
		rom[ 2015 ] =    -77;
		rom[ 2016 ] =    -19;
		rom[ 2017 ] =   -238;
		rom[ 2018 ] =      4;
		rom[ 2019 ] =   -202;
		rom[ 2020 ] =   -487;
		rom[ 2021 ] =    -74;
		rom[ 2022 ] =    -32;
		rom[ 2023 ] =    212;
		rom[ 2024 ] =    273;
		rom[ 2025 ] =    -56;
		rom[ 2026 ] =    -72;
		rom[ 2027 ] =   -172;
		rom[ 2028 ] =    -55;
		rom[ 2029 ] =    -45;
		rom[ 2030 ] =   -503;
		rom[ 2031 ] =    195;
		rom[ 2032 ] =    130;
		rom[ 2033 ] =     17;
		rom[ 2034 ] =   -251;
		rom[ 2035 ] =    -11;
		rom[ 2036 ] =   -280;
		rom[ 2037 ] =    424;
		rom[ 2038 ] =     64;
		rom[ 2039 ] =    -40;
		rom[ 2040 ] =    -36;
		rom[ 2041 ] =   -261;
		rom[ 2042 ] =    159;
		rom[ 2043 ] =   -163;
		rom[ 2044 ] =    206;
		rom[ 2045 ] =    189;
		rom[ 2046 ] =    254;
		rom[ 2047 ] =   -265;
		rom[ 2048 ] =    112;
		rom[ 2049 ] =      1;
		rom[ 2050 ] =    -17;
		rom[ 2051 ] =    193;
		rom[ 2052 ] =     51;
		rom[ 2053 ] =    188;
		rom[ 2054 ] =    813;
		rom[ 2055 ] =     68;
		rom[ 2056 ] =      8;
		rom[ 2057 ] =     91;
		rom[ 2058 ] =    -56;
		rom[ 2059 ] =    -31;
		rom[ 2060 ] =    -54;
		rom[ 2061 ] =    200;
		rom[ 2062 ] =     83;
		rom[ 2063 ] =    -68;
		rom[ 2064 ] =   -693;
		rom[ 2065 ] =   -464;
		rom[ 2066 ] =   -318;
		rom[ 2067 ] =    -63;
		rom[ 2068 ] =   -270;
		rom[ 2069 ] =     34;
		rom[ 2070 ] =    145;
		rom[ 2071 ] =   -159;
		rom[ 2072 ] =    -40;
		rom[ 2073 ] =    -94;
		rom[ 2074 ] =     12;
		rom[ 2075 ] =     53;
		rom[ 2076 ] =     60;
		rom[ 2077 ] =   -246;
		rom[ 2078 ] =    212;
		rom[ 2079 ] =    101;
		rom[ 2080 ] =    -49;
		rom[ 2081 ] =   -404;
		rom[ 2082 ] =    481;
		rom[ 2083 ] =    -77;
		rom[ 2084 ] =   -116;
		rom[ 2085 ] =     53;
		rom[ 2086 ] =   -477;
		rom[ 2087 ] =    -15;
		rom[ 2088 ] =    127;
		rom[ 2089 ] =    103;
		rom[ 2090 ] =   -115;
		rom[ 2091 ] =    149;
		rom[ 2092 ] =   -296;
		rom[ 2093 ] =   -170;
		rom[ 2094 ] =    195;
		rom[ 2095 ] =    269;
		rom[ 2096 ] =     56;
		rom[ 2097 ] =   -113;
		rom[ 2098 ] =    -65;
		rom[ 2099 ] =    303;
		rom[ 2100 ] =     -3;
		rom[ 2101 ] =     73;
		rom[ 2102 ] =    -10;
		rom[ 2103 ] =    -37;
		rom[ 2104 ] =    201;
		rom[ 2105 ] =   -125;
		rom[ 2106 ] =    410;
		rom[ 2107 ] =     13;
		rom[ 2108 ] =    145;
		rom[ 2109 ] =      1;
		rom[ 2110 ] =    103;
		rom[ 2111 ] =    -21;
		rom[ 2112 ] =      6;
		rom[ 2113 ] =    -66;
		rom[ 2114 ] =   -121;
		rom[ 2115 ] =     -6;
		rom[ 2116 ] =   -221;
		rom[ 2117 ] =   -271;
		rom[ 2118 ] =    114;
		rom[ 2119 ] =    118;
		rom[ 2120 ] =    -83;
		rom[ 2121 ] =     50;
		rom[ 2122 ] =    177;
		rom[ 2123 ] =    762;
		rom[ 2124 ] =    130;
		rom[ 2125 ] =     57;
		rom[ 2126 ] =    -25;
		rom[ 2127 ] =    -22;
		rom[ 2128 ] =     68;
		rom[ 2129 ] =    106;
		rom[ 2130 ] =   -109;
		rom[ 2131 ] =    -69;
		rom[ 2132 ] =     24;
		rom[ 2133 ] =    -11;
		rom[ 2134 ] =   -179;
		rom[ 2135 ] =    211;
		rom[ 2136 ] =     33;
		rom[ 2137 ] =   -216;
		rom[ 2138 ] =    215;
		rom[ 2139 ] =    -51;
		rom[ 2140 ] =     47;
		rom[ 2141 ] =    -97;
		rom[ 2142 ] =   -252;
		rom[ 2143 ] =     -7;
		rom[ 2144 ] =    144;
		rom[ 2145 ] =    -75;
		rom[ 2146 ] =   -157;
		rom[ 2147 ] =    408;
		rom[ 2148 ] =    345;
		rom[ 2149 ] =    164;
		rom[ 2150 ] =    241;
		rom[ 2151 ] =    612;
		rom[ 2152 ] =      2;
		rom[ 2153 ] =   -136;
		rom[ 2154 ] =     38;
		rom[ 2155 ] =    176;
		rom[ 2156 ] =   -276;
		rom[ 2157 ] =  -1276;
		rom[ 2158 ] =    121;
		rom[ 2159 ] =     43;
		rom[ 2160 ] =   -118;
		rom[ 2161 ] =    -23;
		rom[ 2162 ] =    116;
		rom[ 2163 ] =   -118;
		rom[ 2164 ] =    102;
		rom[ 2165 ] =     49;
		rom[ 2166 ] =   -174;
		rom[ 2167 ] =     42;
		rom[ 2168 ] =   -283;
		rom[ 2169 ] =    -19;
		rom[ 2170 ] =    -57;
		rom[ 2171 ] =    -62;
		rom[ 2172 ] =    -41;
		rom[ 2173 ] =   -208;
		rom[ 2174 ] =    125;
		rom[ 2175 ] =    -45;
		rom[ 2176 ] =    -25;
		rom[ 2177 ] =    321;
		rom[ 2178 ] =    -41;
		rom[ 2179 ] =    127;
		rom[ 2180 ] =    164;
		rom[ 2181 ] =     66;
		rom[ 2182 ] =   -186;
		rom[ 2183 ] =    -74;
		rom[ 2184 ] =    -57;
		rom[ 2185 ] =   -158;
		rom[ 2186 ] =    129;
		rom[ 2187 ] =    -44;
		rom[ 2188 ] =     49;
		rom[ 2189 ] =    289;
		rom[ 2190 ] =   2176;
		rom[ 2191 ] =    -60;
		rom[ 2192 ] =     -9;
		rom[ 2193 ] =    204;
		rom[ 2194 ] =   -195;
		rom[ 2195 ] =   -374;
		rom[ 2196 ] =    155;
		rom[ 2197 ] =    -63;
		rom[ 2198 ] =    -63;
		rom[ 2199 ] =   -235;
		rom[ 2200 ] =    -24;
		rom[ 2201 ] =   -286;
		rom[ 2202 ] =   -102;
		rom[ 2203 ] =     70;
		rom[ 2204 ] =   -181;
		rom[ 2205 ] =    180;
		rom[ 2206 ] =     65;
		rom[ 2207 ] =   -379;
		rom[ 2208 ] =    290;
		rom[ 2209 ] =    236;
		rom[ 2210 ] =    -67;
		rom[ 2211 ] =     98;
		rom[ 2212 ] =     51;
		rom[ 2213 ] =   -222;
		rom[ 2214 ] =    -54;
		rom[ 2215 ] =     25;
		rom[ 2216 ] =    118;
		rom[ 2217 ] =    -90;
		rom[ 2218 ] =     21;
		rom[ 2219 ] =    352;
		rom[ 2220 ] =    -35;
		rom[ 2221 ] =     27;
		rom[ 2222 ] =    -26;
		rom[ 2223 ] =     36;
		rom[ 2224 ] =     13;
		rom[ 2225 ] =    169;
		rom[ 2226 ] =    -27;
		rom[ 2227 ] =    125;
		rom[ 2228 ] =    -30;
		rom[ 2229 ] =    364;
		rom[ 2230 ] =     29;
		rom[ 2231 ] =    -74;
		rom[ 2232 ] =   -105;
		rom[ 2233 ] =    447;
		rom[ 2234 ] =    -46;
		rom[ 2235 ] =   -235;
		rom[ 2236 ] =    420;
		rom[ 2237 ] =    110;
		rom[ 2238 ] =    -55;
		rom[ 2239 ] =  -1317;
		rom[ 2240 ] =    837;
		rom[ 2241 ] =   -288;
		rom[ 2242 ] =    154;
		rom[ 2243 ] =   -287;
		rom[ 2244 ] =    258;
		rom[ 2245 ] =    149;
		rom[ 2246 ] =     16;
		rom[ 2247 ] =   -201;
		rom[ 2248 ] =   -293;
		rom[ 2249 ] =   -155;
		rom[ 2250 ] =    -12;
		rom[ 2251 ] =     79;
		rom[ 2252 ] =     46;
		rom[ 2253 ] =   -137;
		rom[ 2254 ] =    376;
		rom[ 2255 ] =     15;
		rom[ 2256 ] =     52;
		rom[ 2257 ] =   -586;
		rom[ 2258 ] =   -396;
		rom[ 2259 ] =    -36;
		rom[ 2260 ] =     65;
		rom[ 2261 ] =    288;
		rom[ 2262 ] =   -155;
		rom[ 2263 ] =   2113;
		rom[ 2264 ] =   -134;
		rom[ 2265 ] =   -148;
		rom[ 2266 ] =     27;
		rom[ 2267 ] =    -66;
		rom[ 2268 ] =     34;
		rom[ 2269 ] =   -563;
		rom[ 2270 ] =    724;
		rom[ 2271 ] =     32;
		rom[ 2272 ] =    449;
		rom[ 2273 ] =   -124;
		rom[ 2274 ] =    -94;
		rom[ 2275 ] =    -12;
		rom[ 2276 ] =   -136;
		rom[ 2277 ] =     54;
		rom[ 2278 ] =     60;
		rom[ 2279 ] =    -54;
		rom[ 2280 ] =    -66;
		rom[ 2281 ] =   -118;
		rom[ 2282 ] =   -415;
		rom[ 2283 ] =    154;
		rom[ 2284 ] =  -1169;
		rom[ 2285 ] =    629;
		rom[ 2286 ] =      0;
		rom[ 2287 ] =    -84;
		rom[ 2288 ] =    153;
		rom[ 2289 ] =    234;
		rom[ 2290 ] =     20;
		rom[ 2291 ] =   -223;
		rom[ 2292 ] =    103;
		rom[ 2293 ] =     99;
		rom[ 2294 ] =    147;
		rom[ 2295 ] =   -409;
		rom[ 2296 ] =    345;
		rom[ 2297 ] =     65;
		rom[ 2298 ] =    138;
		rom[ 2299 ] =   -253;
		rom[ 2300 ] =    286;
		rom[ 2301 ] =   -114;
		rom[ 2302 ] =    -52;
		rom[ 2303 ] =     88;
		rom[ 2304 ] =    411;
		rom[ 2305 ] =    106;
		rom[ 2306 ] =    116;
		rom[ 2307 ] =    158;
		rom[ 2308 ] =   -190;
		rom[ 2309 ] =   -175;
		rom[ 2310 ] =     15;
		rom[ 2311 ] =    173;
		rom[ 2312 ] =     80;
		rom[ 2313 ] =      3;
		rom[ 2314 ] =    -17;
		rom[ 2315 ] =     69;
		rom[ 2316 ] =    147;
		rom[ 2317 ] =   -290;
		rom[ 2318 ] =   -258;
		rom[ 2319 ] =    121;
		rom[ 2320 ] =    155;
		rom[ 2321 ] =   -136;
		rom[ 2322 ] =   -129;
		rom[ 2323 ] =      4;
		rom[ 2324 ] =   -293;
		rom[ 2325 ] =   -332;
		rom[ 2326 ] =     18;
		rom[ 2327 ] =   -172;
		rom[ 2328 ] =   -268;
		rom[ 2329 ] =     74;
		rom[ 2330 ] =   -211;
		rom[ 2331 ] =   -193;
		rom[ 2332 ] =     71;
		rom[ 2333 ] =   -103;
		rom[ 2334 ] =   -166;
		rom[ 2335 ] =   -154;
		rom[ 2336 ] =    -54;
		rom[ 2337 ] =      0;
		rom[ 2338 ] =    -46;
		rom[ 2339 ] =    152;
		rom[ 2340 ] =     13;
		rom[ 2341 ] =    -92;
		rom[ 2342 ] =     95;
		rom[ 2343 ] =    -57;
		rom[ 2344 ] =     30;
		rom[ 2345 ] =    -47;
		rom[ 2346 ] =    215;
		rom[ 2347 ] =    215;
		rom[ 2348 ] =    -48;
		rom[ 2349 ] =    392;
		rom[ 2350 ] =    -65;
		rom[ 2351 ] =    142;
		rom[ 2352 ] =    142;
		rom[ 2353 ] =     66;
		rom[ 2354 ] =   -181;
		rom[ 2355 ] =    -22;
		rom[ 2356 ] =   -269;
		rom[ 2357 ] =   -300;
		rom[ 2358 ] =     67;
		rom[ 2359 ] =    -37;
		rom[ 2360 ] =     24;
		rom[ 2361 ] =     -3;
		rom[ 2362 ] =    841;
		rom[ 2363 ] =    -69;
		rom[ 2364 ] =    -78;
		rom[ 2365 ] =   -106;
		rom[ 2366 ] =    -89;
		rom[ 2367 ] =    -98;
		rom[ 2368 ] =    193;
		rom[ 2369 ] =   -188;
		rom[ 2370 ] =    108;
		rom[ 2371 ] =   -199;
		rom[ 2372 ] =    -76;
		rom[ 2373 ] =     51;
		rom[ 2374 ] =     -4;
		rom[ 2375 ] =   -201;
		rom[ 2376 ] =    -71;
		rom[ 2377 ] =    -60;
		rom[ 2378 ] =   -938;
		rom[ 2379 ] =   -520;
		rom[ 2380 ] =     42;
		rom[ 2381 ] =     28;
		rom[ 2382 ] =   1188;
		rom[ 2383 ] =   -975;
		rom[ 2384 ] =    255;
		rom[ 2385 ] =     19;
		rom[ 2386 ] =   -113;
		rom[ 2387 ] =    -69;
		rom[ 2388 ] =   -203;
		rom[ 2389 ] =   -306;
		rom[ 2390 ] =    131;
		rom[ 2391 ] =   -386;
		rom[ 2392 ] =    -63;
		rom[ 2393 ] =    -16;
		rom[ 2394 ] =     12;
		rom[ 2395 ] =    -41;
		rom[ 2396 ] =   -158;
		rom[ 2397 ] =    141;
		rom[ 2398 ] =    -19;
		rom[ 2399 ] =      2;
		rom[ 2400 ] =    144;
		rom[ 2401 ] =    -96;
		rom[ 2402 ] =     -7;
		rom[ 2403 ] =    -68;
		rom[ 2404 ] =   2705;
		rom[ 2405 ] =    449;
		rom[ 2406 ] =     55;
		rom[ 2407 ] =    -93;
		rom[ 2408 ] =   -335;
		rom[ 2409 ] =   -215;
		rom[ 2410 ] =   -103;
		rom[ 2411 ] =   -179;
		rom[ 2412 ] =    -74;
		rom[ 2413 ] =     96;
		rom[ 2414 ] =    140;
		rom[ 2415 ] =    105;
		rom[ 2416 ] =   -108;
		rom[ 2417 ] =    249;
		rom[ 2418 ] =    592;
		rom[ 2419 ] =    218;
		rom[ 2420 ] =     46;
		rom[ 2421 ] =     -9;
		rom[ 2422 ] =   -121;
		rom[ 2423 ] =    111;
		rom[ 2424 ] =    -14;
		rom[ 2425 ] =    -51;
		rom[ 2426 ] =   -363;
		rom[ 2427 ] =    -78;
		rom[ 2428 ] =    -68;
		rom[ 2429 ] =     52;
		rom[ 2430 ] =    -55;
		rom[ 2431 ] =     77;
		rom[ 2432 ] =    -26;
		rom[ 2433 ] =    -99;
		rom[ 2434 ] =   -121;
		rom[ 2435 ] =     20;
		rom[ 2436 ] =    -23;
		rom[ 2437 ] =     68;
		rom[ 2438 ] =    156;
		rom[ 2439 ] =   -233;
		rom[ 2440 ] =   -220;
		rom[ 2441 ] =    -10;
		rom[ 2442 ] =   1217;
		rom[ 2443 ] =   -364;
		rom[ 2444 ] =   -230;
		rom[ 2445 ] =    151;
		rom[ 2446 ] =    -34;
		rom[ 2447 ] =     -9;
		rom[ 2448 ] =   -293;
		rom[ 2449 ] =     21;
		rom[ 2450 ] =    -25;
		rom[ 2451 ] =     63;
		rom[ 2452 ] =    106;
		rom[ 2453 ] =    -49;
		rom[ 2454 ] =   -277;
		rom[ 2455 ] =    -60;
		rom[ 2456 ] =    102;
		rom[ 2457 ] =     77;
		rom[ 2458 ] =    -87;
		rom[ 2459 ] =     38;
		rom[ 2460 ] =    940;
		rom[ 2461 ] =   -155;
		rom[ 2462 ] =    -55;
		rom[ 2463 ] =    148;
		rom[ 2464 ] =     27;
		rom[ 2465 ] =    395;
		rom[ 2466 ] =   -146;
		rom[ 2467 ] =     44;
		rom[ 2468 ] =    324;
		rom[ 2469 ] =    134;
		rom[ 2470 ] =   -113;
		rom[ 2471 ] =    -16;
		rom[ 2472 ] =     30;
		rom[ 2473 ] =    459;
		rom[ 2474 ] =   -486;
		rom[ 2475 ] =   -170;
		rom[ 2476 ] =   -114;
		rom[ 2477 ] =   -512;
		rom[ 2478 ] =    969;
		rom[ 2479 ] =   -120;
		rom[ 2480 ] =    154;
		rom[ 2481 ] =    295;
		rom[ 2482 ] =     40;
		rom[ 2483 ] =    213;
		rom[ 2484 ] =   -179;
		rom[ 2485 ] =   -157;
		rom[ 2486 ] =   -404;
		rom[ 2487 ] =   -499;
		rom[ 2488 ] =   -490;
		rom[ 2489 ] =    126;
		rom[ 2490 ] =     44;
		rom[ 2491 ] =    232;
		rom[ 2492 ] =      4;
		rom[ 2493 ] =   -115;
		rom[ 2494 ] =   -655;
		rom[ 2495 ] =     20;
		rom[ 2496 ] =    192;
		rom[ 2497 ] =     99;
		rom[ 2498 ] =    287;
		rom[ 2499 ] =     40;
		rom[ 2500 ] =   -230;
		rom[ 2501 ] =    449;
		rom[ 2502 ] =     85;
		rom[ 2503 ] =    143;
		rom[ 2504 ] =    163;
		rom[ 2505 ] =    -19;
		rom[ 2506 ] =      9;
		rom[ 2507 ] =    103;
		rom[ 2508 ] =   -131;
		rom[ 2509 ] =    308;
		rom[ 2510 ] =    -75;
		rom[ 2511 ] =    -52;
		rom[ 2512 ] =   -108;
		rom[ 2513 ] =     90;
		rom[ 2514 ] =    600;
		rom[ 2515 ] =     14;
		rom[ 2516 ] =     38;
		rom[ 2517 ] =    -35;
		rom[ 2518 ] =   -160;
		rom[ 2519 ] =    101;
		rom[ 2520 ] =   -143;
		rom[ 2521 ] =    -75;
		rom[ 2522 ] =    -55;
		rom[ 2523 ] =     25;
		rom[ 2524 ] =    -75;
		rom[ 2525 ] =     58;
		rom[ 2526 ] =   -133;
		rom[ 2527 ] =    -10;
		rom[ 2528 ] =     -3;
		rom[ 2529 ] =    194;
		rom[ 2530 ] =    -28;
		rom[ 2531 ] =   -176;
		rom[ 2532 ] =     84;
		rom[ 2533 ] =    -91;
		rom[ 2534 ] =    204;
		rom[ 2535 ] =    253;
		rom[ 2536 ] =   -171;
		rom[ 2537 ] =    -13;
		rom[ 2538 ] =     99;
		rom[ 2539 ] =    -70;
		rom[ 2540 ] =    -16;
		rom[ 2541 ] =    -58;
		rom[ 2542 ] =    -37;
		rom[ 2543 ] =   -506;
		rom[ 2544 ] =   -336;
		rom[ 2545 ] =    268;
		rom[ 2546 ] =   -129;
		rom[ 2547 ] =   -326;
		rom[ 2548 ] =    -77;
		rom[ 2549 ] =    -20;
		rom[ 2550 ] =    -50;
		rom[ 2551 ] =      5;
		rom[ 2552 ] =    121;
		rom[ 2553 ] =    115;
		rom[ 2554 ] =    124;
		rom[ 2555 ] =    -70;
		rom[ 2556 ] =   -344;
		rom[ 2557 ] =     30;
		rom[ 2558 ] =    231;
		rom[ 2559 ] =    -21;
		rom[ 2560 ] =    -61;
		rom[ 2561 ] =    224;
		rom[ 2562 ] =    -80;
		rom[ 2563 ] =   -275;
		rom[ 2564 ] =    -58;
		rom[ 2565 ] =    122;
		rom[ 2566 ] =    212;
		rom[ 2567 ] =    168;
		rom[ 2568 ] =   -526;
		rom[ 2569 ] =      9;
		rom[ 2570 ] =     31;
		rom[ 2571 ] =    186;
		rom[ 2572 ] =   -322;
		rom[ 2573 ] =     32;
		rom[ 2574 ] =    -55;
		rom[ 2575 ] =    118;
		rom[ 2576 ] =   -112;
		rom[ 2577 ] =   -298;
		rom[ 2578 ] =    -57;
		rom[ 2579 ] =    177;
		rom[ 2580 ] =    120;
		rom[ 2581 ] =   -130;
		rom[ 2582 ] =    155;
		rom[ 2583 ] =    -91;
		rom[ 2584 ] =    241;
		rom[ 2585 ] =    127;
		rom[ 2586 ] =    153;
		rom[ 2587 ] =    -85;
		rom[ 2588 ] =   -104;
		rom[ 2589 ] =    -29;
		rom[ 2590 ] =   -208;
		rom[ 2591 ] =    -84;
		rom[ 2592 ] =     43;
		rom[ 2593 ] =    130;
		rom[ 2594 ] =    -97;
		rom[ 2595 ] =    -24;
		rom[ 2596 ] =     97;
		rom[ 2597 ] =    114;
		rom[ 2598 ] =     59;
		rom[ 2599 ] =    445;
		rom[ 2600 ] =    -57;
		rom[ 2601 ] =     16;
		rom[ 2602 ] =    -20;
		rom[ 2603 ] =   -348;
		rom[ 2604 ] =      8;
		rom[ 2605 ] =   1490;
		rom[ 2606 ] =    904;
		rom[ 2607 ] =    -66;
		rom[ 2608 ] =   -197;
		rom[ 2609 ] =     71;
		rom[ 2610 ] =   -140;
		rom[ 2611 ] =    -18;
		rom[ 2612 ] =    528;
		rom[ 2613 ] =    124;
		rom[ 2614 ] =    180;
		rom[ 2615 ] =     12;
		rom[ 2616 ] =   -107;
		rom[ 2617 ] =   -114;
		rom[ 2618 ] =     48;
		rom[ 2619 ] =      6;
		rom[ 2620 ] =    -14;
		rom[ 2621 ] =   -129;
		rom[ 2622 ] =   -131;
		rom[ 2623 ] =    636;
		rom[ 2624 ] =    360;
		rom[ 2625 ] =     -6;
		rom[ 2626 ] =     38;
		rom[ 2627 ] =    152;
		rom[ 2628 ] =    328;
		rom[ 2629 ] =     -3;
		rom[ 2630 ] =    -20;
		rom[ 2631 ] =    489;
		rom[ 2632 ] =    -18;
		rom[ 2633 ] =   -121;
		rom[ 2634 ] =    109;
		rom[ 2635 ] =    181;
		rom[ 2636 ] =    -99;
		rom[ 2637 ] =     80;
		rom[ 2638 ] =     22;
		rom[ 2639 ] =   -950;
		rom[ 2640 ] =   -104;
		rom[ 2641 ] =    -26;
		rom[ 2642 ] =     16;
		rom[ 2643 ] =   -146;
		rom[ 2644 ] =    -58;
		rom[ 2645 ] =   -517;
		rom[ 2646 ] =    281;
		rom[ 2647 ] =    351;
		rom[ 2648 ] =     63;
		rom[ 2649 ] =    332;
		rom[ 2650 ] =     75;
		rom[ 2651 ] =   -353;
		rom[ 2652 ] =    296;
		rom[ 2653 ] =   -320;
		rom[ 2654 ] =    396;
		rom[ 2655 ] =   -163;
		rom[ 2656 ] =    -39;
		rom[ 2657 ] =      1;
		rom[ 2658 ] =     49;
		rom[ 2659 ] =    -85;
		rom[ 2660 ] =    237;
		rom[ 2661 ] =      0;
		rom[ 2662 ] =    -70;
		rom[ 2663 ] =    125;
		rom[ 2664 ] =     -3;
		rom[ 2665 ] =    360;
		rom[ 2666 ] =   -159;
		rom[ 2667 ] =    328;
		rom[ 2668 ] =    161;
		rom[ 2669 ] =     84;
		rom[ 2670 ] =   -274;
		rom[ 2671 ] =    191;
		rom[ 2672 ] =    321;
		rom[ 2673 ] =    271;
		rom[ 2674 ] =    123;
		rom[ 2675 ] =     70;
		rom[ 2676 ] =     82;
		rom[ 2677 ] =    135;
		rom[ 2678 ] =    -60;
		rom[ 2679 ] =    -42;
		rom[ 2680 ] =   -117;
		rom[ 2681 ] =    -19;
		rom[ 2682 ] =   1318;
		rom[ 2683 ] =    -69;
		rom[ 2684 ] =    -30;
		rom[ 2685 ] =   -122;
		rom[ 2686 ] =    -46;
		rom[ 2687 ] =     19;
		rom[ 2688 ] =     20;
		rom[ 2689 ] =    792;
		rom[ 2690 ] =     22;
		rom[ 2691 ] =   -279;
		rom[ 2692 ] =   -143;
		rom[ 2693 ] =     20;
		rom[ 2694 ] =    390;
		rom[ 2695 ] =   -257;
		rom[ 2696 ] =   -697;
		rom[ 2697 ] =     43;
		rom[ 2698 ] =   -170;
		rom[ 2699 ] =    520;
		rom[ 2700 ] =    338;
		rom[ 2701 ] =    349;
		rom[ 2702 ] =    227;
		rom[ 2703 ] =     18;
		rom[ 2704 ] =     53;
		rom[ 2705 ] =    237;
		rom[ 2706 ] =    -93;
		rom[ 2707 ] =    197;
		rom[ 2708 ] =    105;
		rom[ 2709 ] =     28;
		rom[ 2710 ] =   -141;
		rom[ 2711 ] =    120;
		rom[ 2712 ] =     -9;
		rom[ 2713 ] =   -392;
		rom[ 2714 ] =     68;
		rom[ 2715 ] =    106;
		rom[ 2716 ] =      1;
		rom[ 2717 ] =    -27;
		rom[ 2718 ] =     77;
		rom[ 2719 ] =      0;
		rom[ 2720 ] =   -312;
		rom[ 2721 ] =    205;
		rom[ 2722 ] =    -11;
		rom[ 2723 ] =     66;
		rom[ 2724 ] =    154;
		rom[ 2725 ] =    -50;
		rom[ 2726 ] =    237;
		rom[ 2727 ] =     19;
		rom[ 2728 ] =    187;
		rom[ 2729 ] =     87;
		rom[ 2730 ] =    642;
		rom[ 2731 ] =    -42;
		rom[ 2732 ] =      9;
		rom[ 2733 ] =    -95;
		rom[ 2734 ] =    -28;
		rom[ 2735 ] =   -140;
		rom[ 2736 ] =    -86;
		rom[ 2737 ] =      8;
		rom[ 2738 ] =    -17;
		rom[ 2739 ] =    -58;
		rom[ 2740 ] =    -33;
		rom[ 2741 ] =    -38;
		rom[ 2742 ] =   -155;
		rom[ 2743 ] =     19;
		rom[ 2744 ] =    -18;
		rom[ 2745 ] =     21;
		rom[ 2746 ] =    -39;
		rom[ 2747 ] =    184;
		rom[ 2748 ] =     58;
		rom[ 2749 ] =    670;
		rom[ 2750 ] =     10;
		rom[ 2751 ] =    -15;
		rom[ 2752 ] =   -103;
		rom[ 2753 ] =    -79;
		rom[ 2754 ] =     59;
		rom[ 2755 ] =    211;
		rom[ 2756 ] =   -155;
		rom[ 2757 ] =   -121;
		rom[ 2758 ] =   -160;
		rom[ 2759 ] =   -119;
		rom[ 2760 ] =   -342;
		rom[ 2761 ] =   1720;
		rom[ 2762 ] =    245;
		rom[ 2763 ] =    -77;
		rom[ 2764 ] =    -24;
		rom[ 2765 ] =   -238;
		rom[ 2766 ] =    -50;
		rom[ 2767 ] =    190;
		rom[ 2768 ] =      4;
		rom[ 2769 ] =   -363;
		rom[ 2770 ] =    -94;
		rom[ 2771 ] =    176;
		rom[ 2772 ] =      0;
		rom[ 2773 ] =     36;
		rom[ 2774 ] =    -72;
		rom[ 2775 ] =     25;
		rom[ 2776 ] =     93;
		rom[ 2777 ] =    -88;
		rom[ 2778 ] =    252;
		rom[ 2779 ] =   -319;
		rom[ 2780 ] =     46;
		rom[ 2781 ] =   -104;
		rom[ 2782 ] =   -155;
		rom[ 2783 ] =     40;
		rom[ 2784 ] =    -56;
		rom[ 2785 ] =     34;
		rom[ 2786 ] =   -292;
		rom[ 2787 ] =     40;
		rom[ 2788 ] =    450;
		rom[ 2789 ] =    144;
		rom[ 2790 ] =   -457;
		rom[ 2791 ] =   -465;
		rom[ 2792 ] =     68;
		rom[ 2793 ] =    -32;
		rom[ 2794 ] =   -135;
		rom[ 2795 ] =     51;
		rom[ 2796 ] =   -172;
		rom[ 2797 ] =    103;
		rom[ 2798 ] =    -99;
		rom[ 2799 ] =    -50;
		rom[ 2800 ] =   -466;
		rom[ 2801 ] =   -347;
		rom[ 2802 ] =   -100;
		rom[ 2803 ] =    -36;
		rom[ 2804 ] =     45;
		rom[ 2805 ] =   -120;
		rom[ 2806 ] =     26;
		rom[ 2807 ] =     57;
		rom[ 2808 ] =    -54;
		rom[ 2809 ] =   1164;
		rom[ 2810 ] =   -971;
		rom[ 2811 ] =   -457;
		rom[ 2812 ] =    523;
		rom[ 2813 ] =   -257;
		rom[ 2814 ] =     71;
		rom[ 2815 ] =      5;
		rom[ 2816 ] =    112;
		rom[ 2817 ] =   -178;
		rom[ 2818 ] =     45;
		rom[ 2819 ] =     85;
		rom[ 2820 ] =    -91;
		rom[ 2821 ] =    133;
		rom[ 2822 ] =     50;
		rom[ 2823 ] =     34;
		rom[ 2824 ] =    153;
		rom[ 2825 ] =    -57;
		rom[ 2826 ] =    233;
		rom[ 2827 ] =     20;
		rom[ 2828 ] =   -100;
		rom[ 2829 ] =    -46;
		rom[ 2830 ] =    141;
		rom[ 2831 ] =     99;
		rom[ 2832 ] =    -32;
		rom[ 2833 ] =    143;
		rom[ 2834 ] =     18;
		rom[ 2835 ] =   -340;
		rom[ 2836 ] =    -57;
		rom[ 2837 ] =      5;
		rom[ 2838 ] =    -68;
		rom[ 2839 ] =   -314;
		rom[ 2840 ] =   -969;
		rom[ 2841 ] =   -411;
		rom[ 2842 ] =      5;
		rom[ 2843 ] =     90;
		rom[ 2844 ] =   -460;
		rom[ 2845 ] =     67;
		rom[ 2846 ] =    278;
		rom[ 2847 ] =     65;
		rom[ 2848 ] =     19;
		rom[ 2849 ] =     27;
		rom[ 2850 ] =     19;
		rom[ 2851 ] =     10;
		rom[ 2852 ] =     11;
		rom[ 2853 ] =   -123;
		rom[ 2854 ] =     58;
		rom[ 2855 ] =   -247;
		rom[ 2856 ] =    -81;
		rom[ 2857 ] =    127;
		rom[ 2858 ] =     74;
		rom[ 2859 ] =      4;
		rom[ 2860 ] =   -150;
		rom[ 2861 ] =     49;
		rom[ 2862 ] =    306;
		rom[ 2863 ] =   -961;
		rom[ 2864 ] =    577;
		rom[ 2865 ] =     25;
		rom[ 2866 ] =   -234;
		rom[ 2867 ] =   -226;
		rom[ 2868 ] =    -88;
		rom[ 2869 ] =    105;
		rom[ 2870 ] =    -53;
		rom[ 2871 ] =      9;
		rom[ 2872 ] =     36;
		rom[ 2873 ] =    -36;
		rom[ 2874 ] =     16;
		rom[ 2875 ] =    102;
		rom[ 2876 ] =    -24;
		rom[ 2877 ] =     17;
		rom[ 2878 ] =   -138;
		rom[ 2879 ] =    182;
		rom[ 2880 ] =   -167;
		rom[ 2881 ] =    161;
		rom[ 2882 ] =   -288;
		rom[ 2883 ] =    146;
		rom[ 2884 ] =   -175;
		rom[ 2885 ] =    -86;
		rom[ 2886 ] =   -644;
		rom[ 2887 ] =     32;
		rom[ 2888 ] =     96;
		rom[ 2889 ] =    305;
		rom[ 2890 ] =     -2;
		rom[ 2891 ] =    -66;
		rom[ 2892 ] =   -135;
		rom[ 2893 ] =    199;
		rom[ 2894 ] =      9;
		rom[ 2895 ] =    185;
		rom[ 2896 ] =    438;
		rom[ 2897 ] =   -165;
		rom[ 2898 ] =    130;
		rom[ 2899 ] =   -235;
		rom[ 2900 ] =     55;
		rom[ 2901 ] =    292;
		rom[ 2902 ] =    -61;
		rom[ 2903 ] =    -41;
		rom[ 2904 ] =     15;
		rom[ 2905 ] =     66;
		rom[ 2906 ] =   -164;
		rom[ 2907 ] =    110;
		rom[ 2908 ] =    214;
		rom[ 2909 ] =    -78;
		rom[ 2910 ] =    -15;
		rom[ 2911 ] =    310;
		rom[ 2912 ] =    -90;
	end
endmodule

module left_tree_rom(
	input 				clk,
	input		[11:0]	addr,
	output reg	[13:0]	q    // x y w h 5bit*4
	);
	reg					[13:0]	rom [4095:0];
	always @(posedge clk) q <= rom[addr];
	initial begin
		rom[ 0    ] =    534;
		rom[ 1    ] =   -477;
		rom[ 2    ] =   -386;
		rom[ 3    ] =   -223;
		rom[ 4    ] =   -199;
		rom[ 5    ] =    142;
		rom[ 6    ] =   -432;
		rom[ 7    ] =   -378;
		rom[ 8    ] =   -219;
		rom[ 9    ] =    318;
		rom[ 10   ] =   -414;
		rom[ 11   ] =   -497;
		rom[ 12   ] =   -142;
		rom[ 13   ] =     68;
		rom[ 14   ] =   -684;
		rom[ 15   ] =   -277;
		rom[ 16   ] =    -90;
		rom[ 17   ] =    237;
		rom[ 18   ] =    296;
		rom[ 19   ] =   -107;
		rom[ 20   ] =    373;
		rom[ 21   ] =    286;
		rom[ 22   ] =    -89;
		rom[ 23   ] =   -155;
		rom[ 24   ] =     99;
		rom[ 25   ] =   -259;
		rom[ 26   ] =   -421;
		rom[ 27   ] =    118;
		rom[ 28   ] =   -167;
		rom[ 29   ] =   -357;
		rom[ 30   ] =   -129;
		rom[ 31   ] =     93;
		rom[ 32   ] =    -77;
		rom[ 33   ] =   -103;
		rom[ 34   ] =    269;
		rom[ 35   ] =   -416;
		rom[ 36   ] =     72;
		rom[ 37   ] =   -259;
		rom[ 38   ] =    -42;
		rom[ 39   ] =    388;
		rom[ 40   ] =    451;
		rom[ 41   ] =    -80;
		rom[ 42   ] =    -25;
		rom[ 43   ] =   -103;
		rom[ 44   ] =     43;
		rom[ 45   ] =    227;
		rom[ 46   ] =    -95;
		rom[ 47   ] =     16;
		rom[ 48   ] =   -447;
		rom[ 49   ] =   -240;
		rom[ 50   ] =    -13;
		rom[ 51   ] =   -468;
		rom[ 52   ] =    295;
		rom[ 53   ] =   -400;
		rom[ 54   ] =   -147;
		rom[ 55   ] =   -373;
		rom[ 56   ] =   -213;
		rom[ 57   ] =    -80;
		rom[ 58   ] =   -111;
		rom[ 59   ] =    381;
		rom[ 60   ] =   -246;
		rom[ 61   ] =   -626;
		rom[ 62   ] =     44;
		rom[ 63   ] =    124;
		rom[ 64   ] =     45;
		rom[ 65   ] =   -501;
		rom[ 66   ] =    253;
		rom[ 67   ] =   -660;
		rom[ 68   ] =    368;
		rom[ 69   ] =   -126;
		rom[ 70   ] =   -596;
		rom[ 71   ] =   -216;
		rom[ 72   ] =   -369;
		rom[ 73   ] =     46;
		rom[ 74   ] =     17;
		rom[ 75   ] =    100;
		rom[ 76   ] =     37;
		rom[ 77   ] =     63;
		rom[ 78   ] =   -193;
		rom[ 79   ] =    -93;
		rom[ 80   ] =   -594;
		rom[ 81   ] =    108;
		rom[ 82   ] =    284;
		rom[ 83   ] =   -851;
		rom[ 84   ] =   -311;
		rom[ 85   ] =   -123;
		rom[ 86   ] =   -276;
		rom[ 87   ] =   -307;
		rom[ 88   ] =   -112;
		rom[ 89   ] =    -47;
		rom[ 90   ] =     77;
		rom[ 91   ] =    319;
		rom[ 92   ] =   -152;
		rom[ 93   ] =     72;
		rom[ 94   ] =    123;
		rom[ 95   ] =     68;
		rom[ 96   ] =   -335;
		rom[ 97   ] =    116;
		rom[ 98   ] =   -443;
		rom[ 99   ] =    -49;
		rom[ 100  ] =   -412;
		rom[ 101  ] =    190;
		rom[ 102  ] =    -68;
		rom[ 103  ] =    -15;
		rom[ 104  ] =    -89;
		rom[ 105  ] =   -268;
		rom[ 106  ] =    211;
		rom[ 107  ] =     52;
		rom[ 108  ] =     52;
		rom[ 109  ] =   -332;
		rom[ 110  ] =   -335;
		rom[ 111  ] =   -269;
		rom[ 112  ] =   -351;
		rom[ 113  ] =     -9;
		rom[ 114  ] =   -255;
		rom[ 115  ] =    370;
		rom[ 116  ] =    -95;
		rom[ 117  ] =   -147;
		rom[ 118  ] =      4;
		rom[ 119  ] =    -20;
		rom[ 120  ] =   -294;
		rom[ 121  ] =     95;
		rom[ 122  ] =     67;
		rom[ 123  ] =    193;
		rom[ 124  ] =     57;
		rom[ 125  ] =   -323;
		rom[ 126  ] =    222;
		rom[ 127  ] =   -355;
		rom[ 128  ] =     16;
		rom[ 129  ] =   -137;
		rom[ 130  ] =    -90;
		rom[ 131  ] =   -150;
		rom[ 132  ] =    -85;
		rom[ 133  ] =    178;
		rom[ 134  ] =    220;
		rom[ 135  ] =     49;
		rom[ 136  ] =   -228;
		rom[ 137  ] =   -322;
		rom[ 138  ] =   -220;
		rom[ 139  ] =   -191;
		rom[ 140  ] =   -323;
		rom[ 141  ] =   -251;
		rom[ 142  ] =    164;
		rom[ 143  ] =    -61;
		rom[ 144  ] =    -87;
		rom[ 145  ] =    281;
		rom[ 146  ] =    402;
		rom[ 147  ] =    -70;
		rom[ 148  ] =   -280;
		rom[ 149  ] =     78;
		rom[ 150  ] =     66;
		rom[ 151  ] =   -315;
		rom[ 152  ] =    104;
		rom[ 153  ] =    -24;
		rom[ 154  ] =   -105;
		rom[ 155  ] =     64;
		rom[ 156  ] =   -240;
		rom[ 157  ] =    318;
		rom[ 158  ] =    -83;
		rom[ 159  ] =     89;
		rom[ 160  ] =     14;
		rom[ 161  ] =   -262;
		rom[ 162  ] =    263;
		rom[ 163  ] =     55;
		rom[ 164  ] =   -408;
		rom[ 165  ] =   -263;
		rom[ 166  ] =   -378;
		rom[ 167  ] =    -61;
		rom[ 168  ] =     74;
		rom[ 169  ] =    -59;
		rom[ 170  ] =   -309;
		rom[ 171  ] =     62;
		rom[ 172  ] =   -350;
		rom[ 173  ] =     54;
		rom[ 174  ] =     83;
		rom[ 175  ] =    -72;
		rom[ 176  ] =   -591;
		rom[ 177  ] =     73;
		rom[ 178  ] =    -69;
		rom[ 179  ] =   -392;
		rom[ 180  ] =     19;
		rom[ 181  ] =     36;
		rom[ 182  ] =   -282;
		rom[ 183  ] =      3;
		rom[ 184  ] =    -88;
		rom[ 185  ] =     51;
		rom[ 186  ] =   -104;
		rom[ 187  ] =   -569;
		rom[ 188  ] =    -73;
		rom[ 189  ] =   -227;
		rom[ 190  ] =   -285;
		rom[ 191  ] =   -258;
		rom[ 192  ] =     66;
		rom[ 193  ] =   -146;
		rom[ 194  ] =   -141;
		rom[ 195  ] =   -329;
		rom[ 196  ] =    446;
		rom[ 197  ] =   -269;
		rom[ 198  ] =    145;
		rom[ 199  ] =    334;
		rom[ 200  ] =   -118;
		rom[ 201  ] =   -106;
		rom[ 202  ] =     92;
		rom[ 203  ] =   -228;
		rom[ 204  ] =     75;
		rom[ 205  ] =   -203;
		rom[ 206  ] =     39;
		rom[ 207  ] =      8;
		rom[ 208  ] =   -100;
		rom[ 209  ] =     22;
		rom[ 210  ] =    141;
		rom[ 211  ] =   -473;
		rom[ 212  ] =   -123;
		rom[ 213  ] =   -115;
		rom[ 214  ] =   -216;
		rom[ 215  ] =     90;
		rom[ 216  ] =     47;
		rom[ 217  ] =   -320;
		rom[ 218  ] =   -208;
		rom[ 219  ] =   -237;
		rom[ 220  ] =    144;
		rom[ 221  ] =    205;
		rom[ 222  ] =   -217;
		rom[ 223  ] =   -103;
		rom[ 224  ] =   -391;
		rom[ 225  ] =    161;
		rom[ 226  ] =    150;
		rom[ 227  ] =    -65;
		rom[ 228  ] =     74;
		rom[ 229  ] =   -101;
		rom[ 230  ] =     53;
		rom[ 231  ] =    112;
		rom[ 232  ] =    240;
		rom[ 233  ] =      2;
		rom[ 234  ] =   -259;
		rom[ 235  ] =    -96;
		rom[ 236  ] =   -206;
		rom[ 237  ] =   -270;
		rom[ 238  ] =     51;
		rom[ 239  ] =    -97;
		rom[ 240  ] =     54;
		rom[ 241  ] =   -262;
		rom[ 242  ] =   -263;
		rom[ 243  ] =    -53;
		rom[ 244  ] =    225;
		rom[ 245  ] =    267;
		rom[ 246  ] =     35;
		rom[ 247  ] =   -425;
		rom[ 248  ] =    204;
		rom[ 249  ] =   -245;
		rom[ 250  ] =     50;
		rom[ 251  ] =   -265;
		rom[ 252  ] =   -315;
		rom[ 253  ] =   -194;
		rom[ 254  ] =    -99;
		rom[ 255  ] =   -183;
		rom[ 256  ] =    141;
		rom[ 257  ] =   -114;
		rom[ 258  ] =   -279;
		rom[ 259  ] =    214;
		rom[ 260  ] =    -65;
		rom[ 261  ] =     80;
		rom[ 262  ] =   -268;
		rom[ 263  ] =     41;
		rom[ 264  ] =   -176;
		rom[ 265  ] =     63;
		rom[ 266  ] =   -129;
		rom[ 267  ] =     10;
		rom[ 268  ] =     36;
		rom[ 269  ] =   -229;
		rom[ 270  ] =   -116;
		rom[ 271  ] =     86;
		rom[ 272  ] =   -202;
		rom[ 273  ] =   -584;
		rom[ 274  ] =    100;
		rom[ 275  ] =      8;
		rom[ 276  ] =   -277;
		rom[ 277  ] =   -481;
		rom[ 278  ] =     37;
		rom[ 279  ] =   -260;
		rom[ 280  ] =     39;
		rom[ 281  ] =   -197;
		rom[ 282  ] =    -29;
		rom[ 283  ] =     17;
		rom[ 284  ] =   -450;
		rom[ 285  ] =    245;
		rom[ 286  ] =    119;
		rom[ 287  ] =    181;
		rom[ 288  ] =   -281;
		rom[ 289  ] =   -279;
		rom[ 290  ] =    -67;
		rom[ 291  ] =    -56;
		rom[ 292  ] =     47;
		rom[ 293  ] =   -237;
		rom[ 294  ] =    502;
		rom[ 295  ] =     54;
		rom[ 296  ] =   -300;
		rom[ 297  ] =   -287;
		rom[ 298  ] =    -43;
		rom[ 299  ] =    211;
		rom[ 300  ] =   -295;
		rom[ 301  ] =   -268;
		rom[ 302  ] =   -279;
		rom[ 303  ] =    108;
		rom[ 304  ] =   -235;
		rom[ 305  ] =   -408;
		rom[ 306  ] =   -169;
		rom[ 307  ] =     49;
		rom[ 308  ] =   -162;
		rom[ 309  ] =    -48;
		rom[ 310  ] =    -27;
		rom[ 311  ] =   -276;
		rom[ 312  ] =     87;
		rom[ 313  ] =    121;
		rom[ 314  ] =    249;
		rom[ 315  ] =   -556;
		rom[ 316  ] =   -164;
		rom[ 317  ] =   -377;
		rom[ 318  ] =    108;
		rom[ 319  ] =      6;
		rom[ 320  ] =     40;
		rom[ 321  ] =   -103;
		rom[ 322  ] =   -510;
		rom[ 323  ] =   -159;
		rom[ 324  ] =    259;
		rom[ 325  ] =   -262;
		rom[ 326  ] =   -291;
		rom[ 327  ] =   -145;
		rom[ 328  ] =     78;
		rom[ 329  ] =   -440;
		rom[ 330  ] =     59;
		rom[ 331  ] =   -311;
		rom[ 332  ] =     83;
		rom[ 333  ] =    -81;
		rom[ 334  ] =    -28;
		rom[ 335  ] =    101;
		rom[ 336  ] =      0;
		rom[ 337  ] =    192;
		rom[ 338  ] =   -212;
		rom[ 339  ] =   -152;
		rom[ 340  ] =     40;
		rom[ 341  ] =      8;
		rom[ 342  ] =   -133;
		rom[ 343  ] =   -136;
		rom[ 344  ] =     51;
		rom[ 345  ] =     11;
		rom[ 346  ] =   -233;
		rom[ 347  ] =     23;
		rom[ 348  ] =     54;
		rom[ 349  ] =    -69;
		rom[ 350  ] =    -26;
		rom[ 351  ] =     16;
		rom[ 352  ] =   -237;
		rom[ 353  ] =     34;
		rom[ 354  ] =     50;
		rom[ 355  ] =   -292;
		rom[ 356  ] =     43;
		rom[ 357  ] =   -121;
		rom[ 358  ] =   -553;
		rom[ 359  ] =     11;
		rom[ 360  ] =     -8;
		rom[ 361  ] =   -337;
		rom[ 362  ] =     94;
		rom[ 363  ] =    -65;
		rom[ 364  ] =    -19;
		rom[ 365  ] =   -201;
		rom[ 366  ] =    435;
		rom[ 367  ] =    198;
		rom[ 368  ] =   -382;
		rom[ 369  ] =   -546;
		rom[ 370  ] =    145;
		rom[ 371  ] =    173;
		rom[ 372  ] =     63;
		rom[ 373  ] =      3;
		rom[ 374  ] =     -2;
		rom[ 375  ] =    115;
		rom[ 376  ] =   -243;
		rom[ 377  ] =   -515;
		rom[ 378  ] =    101;
		rom[ 379  ] =    -63;
		rom[ 380  ] =    -14;
		rom[ 381  ] =     11;
		rom[ 382  ] =   -125;
		rom[ 383  ] =    -76;
		rom[ 384  ] =   -153;
		rom[ 385  ] =     -7;
		rom[ 386  ] =     95;
		rom[ 387  ] =   -255;
		rom[ 388  ] =     36;
		rom[ 389  ] =    -54;
		rom[ 390  ] =   -337;
		rom[ 391  ] =    126;
		rom[ 392  ] =    108;
		rom[ 393  ] =     -7;
		rom[ 394  ] =   -202;
		rom[ 395  ] =   -576;
		rom[ 396  ] =    -65;
		rom[ 397  ] =    -57;
		rom[ 398  ] =    -73;
		rom[ 399  ] =     -8;
		rom[ 400  ] =    152;
		rom[ 401  ] =   -122;
		rom[ 402  ] =     58;
		rom[ 403  ] =    -66;
		rom[ 404  ] =   -153;
		rom[ 405  ] =    181;
		rom[ 406  ] =   -143;
		rom[ 407  ] =   -182;
		rom[ 408  ] =   -285;
		rom[ 409  ] =   -104;
		rom[ 410  ] =    -97;
		rom[ 411  ] =   -179;
		rom[ 412  ] =   -139;
		rom[ 413  ] =    -25;
		rom[ 414  ] =    216;
		rom[ 415  ] =     67;
		rom[ 416  ] =     39;
		rom[ 417  ] =   -509;
		rom[ 418  ] =    -82;
		rom[ 419  ] =    152;
		rom[ 420  ] =      5;
		rom[ 421  ] =   -112;
		rom[ 422  ] =   -228;
		rom[ 423  ] =     54;
		rom[ 424  ] =      3;
		rom[ 425  ] =    257;
		rom[ 426  ] =   -376;
		rom[ 427  ] =   -208;
		rom[ 428  ] =     29;
		rom[ 429  ] =     33;
		rom[ 430  ] =   -301;
		rom[ 431  ] =    161;
		rom[ 432  ] =     47;
		rom[ 433  ] =   -238;
		rom[ 434  ] =      9;
		rom[ 435  ] =     93;
		rom[ 436  ] =     50;
		rom[ 437  ] =   -429;
		rom[ 438  ] =   -787;
		rom[ 439  ] =     54;
		rom[ 440  ] =   -293;
		rom[ 441  ] =    214;
		rom[ 442  ] =    -71;
		rom[ 443  ] =     45;
		rom[ 444  ] =    246;
		rom[ 445  ] =      2;
		rom[ 446  ] =   -136;
		rom[ 447  ] =    210;
		rom[ 448  ] =    -50;
		rom[ 449  ] =     -6;
		rom[ 450  ] =   -347;
		rom[ 451  ] =   -165;
		rom[ 452  ] =    215;
		rom[ 453  ] =     49;
		rom[ 454  ] =   -186;
		rom[ 455  ] =    -92;
		rom[ 456  ] =     14;
		rom[ 457  ] =    120;
		rom[ 458  ] =   -290;
		rom[ 459  ] =    251;
		rom[ 460  ] =    -72;
		rom[ 461  ] =   -163;
		rom[ 462  ] =     95;
		rom[ 463  ] =   -334;
		rom[ 464  ] =   -523;
		rom[ 465  ] =    198;
		rom[ 466  ] =     44;
		rom[ 467  ] =   -384;
		rom[ 468  ] =     73;
		rom[ 469  ] =    354;
		rom[ 470  ] =    -57;
		rom[ 471  ] =   -406;
		rom[ 472  ] =   -305;
		rom[ 473  ] =    -39;
		rom[ 474  ] =     66;
		rom[ 475  ] =    -22;
		rom[ 476  ] =    192;
		rom[ 477  ] =     31;
		rom[ 478  ] =    -93;
		rom[ 479  ] =    -19;
		rom[ 480  ] =    200;
		rom[ 481  ] =   -229;
		rom[ 482  ] =    211;
		rom[ 483  ] =      4;
		rom[ 484  ] =    289;
		rom[ 485  ] =   -147;
		rom[ 486  ] =     -5;
		rom[ 487  ] =   -139;
		rom[ 488  ] =   -313;
		rom[ 489  ] =     37;
		rom[ 490  ] =    -71;
		rom[ 491  ] =    -62;
		rom[ 492  ] =   -219;
		rom[ 493  ] =    177;
		rom[ 494  ] =    -42;
		rom[ 495  ] =    112;
		rom[ 496  ] =   -250;
		rom[ 497  ] =   -231;
		rom[ 498  ] =   -202;
		rom[ 499  ] =    -77;
		rom[ 500  ] =   -230;
		rom[ 501  ] =   -107;
		rom[ 502  ] =    117;
		rom[ 503  ] =    233;
		rom[ 504  ] =   -376;
		rom[ 505  ] =   -268;
		rom[ 506  ] =     74;
		rom[ 507  ] =   -329;
		rom[ 508  ] =   -219;
		rom[ 509  ] =     41;
		rom[ 510  ] =     40;
		rom[ 511  ] =      5;
		rom[ 512  ] =    -42;
		rom[ 513  ] =   -249;
		rom[ 514  ] =    252;
		rom[ 515  ] =    121;
		rom[ 516  ] =   -245;
		rom[ 517  ] =   -134;
		rom[ 518  ] =     43;
		rom[ 519  ] =   -290;
		rom[ 520  ] =     66;
		rom[ 521  ] =     50;
		rom[ 522  ] =    -13;
		rom[ 523  ] =    272;
		rom[ 524  ] =    -47;
		rom[ 525  ] =     -7;
		rom[ 526  ] =    255;
		rom[ 527  ] =     -7;
		rom[ 528  ] =      0;
		rom[ 529  ] =   -391;
		rom[ 530  ] =      8;
		rom[ 531  ] =    196;
		rom[ 532  ] =     41;
		rom[ 533  ] =   -250;
		rom[ 534  ] =    118;
		rom[ 535  ] =     65;
		rom[ 536  ] =   -206;
		rom[ 537  ] =   -336;
		rom[ 538  ] =     51;
		rom[ 539  ] =    249;
		rom[ 540  ] =    -48;
		rom[ 541  ] =   -174;
		rom[ 542  ] =     48;
		rom[ 543  ] =    -60;
		rom[ 544  ] =     63;
		rom[ 545  ] =   -266;
		rom[ 546  ] =    131;
		rom[ 547  ] =    414;
		rom[ 548  ] =    764;
		rom[ 549  ] =    154;
		rom[ 550  ] =   -158;
		rom[ 551  ] =    169;
		rom[ 552  ] =   -287;
		rom[ 553  ] =   -275;
		rom[ 554  ] =    207;
		rom[ 555  ] =     -5;
		rom[ 556  ] =    173;
		rom[ 557  ] =     14;
		rom[ 558  ] =    -33;
		rom[ 559  ] =    -96;
		rom[ 560  ] =   -149;
		rom[ 561  ] =    -77;
		rom[ 562  ] =    151;
		rom[ 563  ] =    248;
		rom[ 564  ] =    233;
		rom[ 565  ] =   -154;
		rom[ 566  ] =     11;
		rom[ 567  ] =   -239;
		rom[ 568  ] =     46;
		rom[ 569  ] =   -330;
		rom[ 570  ] =    -11;
		rom[ 571  ] =     -3;
		rom[ 572  ] =    -68;
		rom[ 573  ] =   -131;
		rom[ 574  ] =    106;
		rom[ 575  ] =    -63;
		rom[ 576  ] =    -57;
		rom[ 577  ] =     16;
		rom[ 578  ] =     48;
		rom[ 579  ] =   -242;
		rom[ 580  ] =     94;
		rom[ 581  ] =    246;
		rom[ 582  ] =   -785;
		rom[ 583  ] =     58;
		rom[ 584  ] =      0;
		rom[ 585  ] =    243;
		rom[ 586  ] =    -25;
		rom[ 587  ] =      2;
		rom[ 588  ] =    165;
		rom[ 589  ] =     -9;
		rom[ 590  ] =    177;
		rom[ 591  ] =   -103;
		rom[ 592  ] =   -165;
		rom[ 593  ] =    250;
		rom[ 594  ] =    -26;
		rom[ 595  ] =    156;
		rom[ 596  ] =   -260;
		rom[ 597  ] =   -105;
		rom[ 598  ] =   -149;
		rom[ 599  ] =   -237;
		rom[ 600  ] =     30;
		rom[ 601  ] =   -148;
		rom[ 602  ] =    -98;
		rom[ 603  ] =    301;
		rom[ 604  ] =   -220;
		rom[ 605  ] =   -191;
		rom[ 606  ] =    235;
		rom[ 607  ] =     68;
		rom[ 608  ] =    -72;
		rom[ 609  ] =   -157;
		rom[ 610  ] =    147;
		rom[ 611  ] =     83;
		rom[ 612  ] =     22;
		rom[ 613  ] =     88;
		rom[ 614  ] =     60;
		rom[ 615  ] =   -190;
		rom[ 616  ] =   -231;
		rom[ 617  ] =    -88;
		rom[ 618  ] =   -239;
		rom[ 619  ] =   -136;
		rom[ 620  ] =    235;
		rom[ 621  ] =   -181;
		rom[ 622  ] =   -222;
		rom[ 623  ] =    -58;
		rom[ 624  ] =    -77;
		rom[ 625  ] =     68;
		rom[ 626  ] =   -302;
		rom[ 627  ] =   -139;
		rom[ 628  ] =    -69;
		rom[ 629  ] =   -233;
		rom[ 630  ] =   -112;
		rom[ 631  ] =      6;
		rom[ 632  ] =    202;
		rom[ 633  ] =    205;
		rom[ 634  ] =    -51;
		rom[ 635  ] =    -11;
		rom[ 636  ] =   -231;
		rom[ 637  ] =     90;
		rom[ 638  ] =    -50;
		rom[ 639  ] =   -358;
		rom[ 640  ] =      0;
		rom[ 641  ] =   -125;
		rom[ 642  ] =   -312;
		rom[ 643  ] =     95;
		rom[ 644  ] =    -75;
		rom[ 645  ] =   -368;
		rom[ 646  ] =   -577;
		rom[ 647  ] =     96;
		rom[ 648  ] =    -75;
		rom[ 649  ] =   -255;
		rom[ 650  ] =     12;
		rom[ 651  ] =     38;
		rom[ 652  ] =     -3;
		rom[ 653  ] =    -36;
		rom[ 654  ] =     -4;
		rom[ 655  ] =   -443;
		rom[ 656  ] =    -61;
		rom[ 657  ] =      1;
		rom[ 658  ] =      9;
		rom[ 659  ] =     19;
		rom[ 660  ] =   -434;
		rom[ 661  ] =    161;
		rom[ 662  ] =    -85;
		rom[ 663  ] =     58;
		rom[ 664  ] =     49;
		rom[ 665  ] =     23;
		rom[ 666  ] =   -446;
		rom[ 667  ] =    -61;
		rom[ 668  ] =    301;
		rom[ 669  ] =     35;
		rom[ 670  ] =   -139;
		rom[ 671  ] =    -55;
		rom[ 672  ] =     16;
		rom[ 673  ] =    175;
		rom[ 674  ] =    445;
		rom[ 675  ] =     78;
		rom[ 676  ] =    -54;
		rom[ 677  ] =   -203;
		rom[ 678  ] =     95;
		rom[ 679  ] =     -3;
		rom[ 680  ] =    310;
		rom[ 681  ] =     -5;
		rom[ 682  ] =   -271;
		rom[ 683  ] =     -8;
		rom[ 684  ] =      9;
		rom[ 685  ] =    -20;
		rom[ 686  ] =   -491;
		rom[ 687  ] =    123;
		rom[ 688  ] =    -50;
		rom[ 689  ] =     50;
		rom[ 690  ] =    -49;
		rom[ 691  ] =    463;
		rom[ 692  ] =    199;
		rom[ 693  ] =     39;
		rom[ 694  ] =    -42;
		rom[ 695  ] =    -26;
		rom[ 696  ] =     -9;
		rom[ 697  ] =    -14;
		rom[ 698  ] =     71;
		rom[ 699  ] =     32;
		rom[ 700  ] =      5;
		rom[ 701  ] =     48;
		rom[ 702  ] =     18;
		rom[ 703  ] =     12;
		rom[ 704  ] =    -69;
		rom[ 705  ] =     13;
		rom[ 706  ] =     97;
		rom[ 707  ] =     39;
		rom[ 708  ] =      6;
		rom[ 709  ] =     41;
		rom[ 710  ] =   -157;
		rom[ 711  ] =   -217;
		rom[ 712  ] =   -208;
		rom[ 713  ] =    -93;
		rom[ 714  ] =   -304;
		rom[ 715  ] =     84;
		rom[ 716  ] =   -130;
		rom[ 717  ] =   -268;
		rom[ 718  ] =   -129;
		rom[ 719  ] =   -254;
		rom[ 720  ] =    -24;
		rom[ 721  ] =     59;
		rom[ 722  ] =    -26;
		rom[ 723  ] =      0;
		rom[ 724  ] =   -167;
		rom[ 725  ] =     72;
		rom[ 726  ] =     39;
		rom[ 727  ] =    -74;
		rom[ 728  ] =    349;
		rom[ 729  ] =    312;
		rom[ 730  ] =   -209;
		rom[ 731  ] =   -312;
		rom[ 732  ] =     30;
		rom[ 733  ] =   -299;
		rom[ 734  ] =   -273;
		rom[ 735  ] =    -92;
		rom[ 736  ] =    125;
		rom[ 737  ] =    150;
		rom[ 738  ] =    -19;
		rom[ 739  ] =     70;
		rom[ 740  ] =     -1;
		rom[ 741  ] =    210;
		rom[ 742  ] =     33;
		rom[ 743  ] =   -232;
		rom[ 744  ] =      2;
		rom[ 745  ] =    455;
		rom[ 746  ] =    146;
		rom[ 747  ] =    -82;
		rom[ 748  ] =     49;
		rom[ 749  ] =     17;
		rom[ 750  ] =    -99;
		rom[ 751  ] =     -6;
		rom[ 752  ] =   -491;
		rom[ 753  ] =   -328;
		rom[ 754  ] =   -103;
		rom[ 755  ] =   -186;
		rom[ 756  ] =    148;
		rom[ 757  ] =    234;
		rom[ 758  ] =   -132;
		rom[ 759  ] =     61;
		rom[ 760  ] =     42;
		rom[ 761  ] =   -349;
		rom[ 762  ] =   -437;
		rom[ 763  ] =    -80;
		rom[ 764  ] =     38;
		rom[ 765  ] =    190;
		rom[ 766  ] =   -104;
		rom[ 767  ] =    208;
		rom[ 768  ] =     84;
		rom[ 769  ] =   -321;
		rom[ 770  ] =    353;
		rom[ 771  ] =     -9;
		rom[ 772  ] =    -47;
		rom[ 773  ] =   -114;
		rom[ 774  ] =    173;
		rom[ 775  ] =     -3;
		rom[ 776  ] =     86;
		rom[ 777  ] =   -271;
		rom[ 778  ] =     37;
		rom[ 779  ] =    -62;
		rom[ 780  ] =     33;
		rom[ 781  ] =   -268;
		rom[ 782  ] =   -387;
		rom[ 783  ] =     35;
		rom[ 784  ] =     73;
		rom[ 785  ] =    -69;
		rom[ 786  ] =     47;
		rom[ 787  ] =     83;
		rom[ 788  ] =     29;
		rom[ 789  ] =   -283;
		rom[ 790  ] =    205;
		rom[ 791  ] =    -67;
		rom[ 792  ] =      4;
		rom[ 793  ] =      3;
		rom[ 794  ] =    -78;
		rom[ 795  ] =   -411;
		rom[ 796  ] =     19;
		rom[ 797  ] =     -1;
		rom[ 798  ] =    -61;
		rom[ 799  ] =    490;
		rom[ 800  ] =    -64;
		rom[ 801  ] =   -177;
		rom[ 802  ] =     46;
		rom[ 803  ] =     -7;
		rom[ 804  ] =     16;
		rom[ 805  ] =      2;
		rom[ 806  ] =     38;
		rom[ 807  ] =     99;
		rom[ 808  ] =   -397;
		rom[ 809  ] =     55;
		rom[ 810  ] =    -12;
		rom[ 811  ] =    -65;
		rom[ 812  ] =    -46;
		rom[ 813  ] =    139;
		rom[ 814  ] =   -177;
		rom[ 815  ] =     75;
		rom[ 816  ] =    236;
		rom[ 817  ] =   -203;
		rom[ 818  ] =     84;
		rom[ 819  ] =   -351;
		rom[ 820  ] =     16;
		rom[ 821  ] =     92;
		rom[ 822  ] =    -39;
		rom[ 823  ] =     34;
		rom[ 824  ] =     27;
		rom[ 825  ] =     -2;
		rom[ 826  ] =      0;
		rom[ 827  ] =   -120;
		rom[ 828  ] =     -2;
		rom[ 829  ] =    -88;
		rom[ 830  ] =    383;
		rom[ 831  ] =   -254;
		rom[ 832  ] =   -147;
		rom[ 833  ] =     -8;
		rom[ 834  ] =    102;
		rom[ 835  ] =     46;
		rom[ 836  ] =    139;
		rom[ 837  ] =    174;
		rom[ 838  ] =   -230;
		rom[ 839  ] =   -144;
		rom[ 840  ] =     92;
		rom[ 841  ] =   -142;
		rom[ 842  ] =   -274;
		rom[ 843  ] =   -183;
		rom[ 844  ] =   -120;
		rom[ 845  ] =     54;
		rom[ 846  ] =    171;
		rom[ 847  ] =   -244;
		rom[ 848  ] =    208;
		rom[ 849  ] =    315;
		rom[ 850  ] =    -78;
		rom[ 851  ] =     54;
		rom[ 852  ] =   -231;
		rom[ 853  ] =     57;
		rom[ 854  ] =   -101;
		rom[ 855  ] =     47;
		rom[ 856  ] =     39;
		rom[ 857  ] =     55;
		rom[ 858  ] =   -378;
		rom[ 859  ] =    -43;
		rom[ 860  ] =      9;
		rom[ 861  ] =     85;
		rom[ 862  ] =      1;
		rom[ 863  ] =    115;
		rom[ 864  ] =     39;
		rom[ 865  ] =   -333;
		rom[ 866  ] =    -62;
		rom[ 867  ] =      7;
		rom[ 868  ] =    -57;
		rom[ 869  ] =     52;
		rom[ 870  ] =    175;
		rom[ 871  ] =     -2;
		rom[ 872  ] =    -51;
		rom[ 873  ] =    121;
		rom[ 874  ] =   -283;
		rom[ 875  ] =    259;
		rom[ 876  ] =    106;
		rom[ 877  ] =     54;
		rom[ 878  ] =   -296;
		rom[ 879  ] =     90;
		rom[ 880  ] =   -393;
		rom[ 881  ] =     51;
		rom[ 882  ] =     -6;
		rom[ 883  ] =     43;
		rom[ 884  ] =   -306;
		rom[ 885  ] =   -279;
		rom[ 886  ] =     71;
		rom[ 887  ] =    -11;
		rom[ 888  ] =    -67;
		rom[ 889  ] =    154;
		rom[ 890  ] =     97;
		rom[ 891  ] =     33;
		rom[ 892  ] =     30;
		rom[ 893  ] =    -87;
		rom[ 894  ] =    -43;
		rom[ 895  ] =    156;
		rom[ 896  ] =   -124;
		rom[ 897  ] =  -1030;
		rom[ 898  ] =   -100;
		rom[ 899  ] =    -22;
		rom[ 900  ] =    293;
		rom[ 901  ] =     -5;
		rom[ 902  ] =      9;
		rom[ 903  ] =    144;
		rom[ 904  ] =    -44;
		rom[ 905  ] =    323;
		rom[ 906  ] =    171;
		rom[ 907  ] =   -105;
		rom[ 908  ] =   -234;
		rom[ 909  ] =      0;
		rom[ 910  ] =    -95;
		rom[ 911  ] =   -108;
		rom[ 912  ] =    -42;
		rom[ 913  ] =     38;
		rom[ 914  ] =    352;
		rom[ 915  ] =    -86;
		rom[ 916  ] =    195;
		rom[ 917  ] =   -177;
		rom[ 918  ] =     -3;
		rom[ 919  ] =    -26;
		rom[ 920  ] =    273;
		rom[ 921  ] =     47;
		rom[ 922  ] =    -56;
		rom[ 923  ] =     65;
		rom[ 924  ] =     -2;
		rom[ 925  ] =    -73;
		rom[ 926  ] =     -9;
		rom[ 927  ] =     84;
		rom[ 928  ] =    -89;
		rom[ 929  ] =   -368;
		rom[ 930  ] =   -302;
		rom[ 931  ] =    566;
		rom[ 932  ] =   -478;
		rom[ 933  ] =   -196;
		rom[ 934  ] =   -161;
		rom[ 935  ] =    218;
		rom[ 936  ] =     -8;
		rom[ 937  ] =    -49;
		rom[ 938  ] =    527;
		rom[ 939  ] =    -29;
		rom[ 940  ] =     -4;
		rom[ 941  ] =    -10;
		rom[ 942  ] =   -170;
		rom[ 943  ] =    -14;
		rom[ 944  ] =    156;
		rom[ 945  ] =   -146;
		rom[ 946  ] =     14;
		rom[ 947  ] =     44;
		rom[ 948  ] =   -171;
		rom[ 949  ] =     75;
		rom[ 950  ] =    -72;
		rom[ 951  ] =    -27;
		rom[ 952  ] =    -13;
		rom[ 953  ] =    115;
		rom[ 954  ] =   -520;
		rom[ 955  ] =     43;
		rom[ 956  ] =     -5;
		rom[ 957  ] =     77;
		rom[ 958  ] =    -79;
		rom[ 959  ] =   -460;
		rom[ 960  ] =    -13;
		rom[ 961  ] =     53;
		rom[ 962  ] =    -51;
		rom[ 963  ] =   -244;
		rom[ 964  ] =    -36;
		rom[ 965  ] =   -279;
		rom[ 966  ] =     26;
		rom[ 967  ] =     15;
		rom[ 968  ] =   -343;
		rom[ 969  ] =     12;
		rom[ 970  ] =   -262;
		rom[ 971  ] =     21;
		rom[ 972  ] =    -37;
		rom[ 973  ] =    168;
		rom[ 974  ] =   -232;
		rom[ 975  ] =   -127;
		rom[ 976  ] =   -108;
		rom[ 977  ] =   -122;
		rom[ 978  ] =    130;
		rom[ 979  ] =    -59;
		rom[ 980  ] =    103;
		rom[ 981  ] =    115;
		rom[ 982  ] =   -217;
		rom[ 983  ] =   -238;
		rom[ 984  ] =   -327;
		rom[ 985  ] =    149;
		rom[ 986  ] =    -13;
		rom[ 987  ] =   -222;
		rom[ 988  ] =    -19;
		rom[ 989  ] =    -63;
		rom[ 990  ] =   -287;
		rom[ 991  ] =   -371;
		rom[ 992  ] =    137;
		rom[ 993  ] =     17;
		rom[ 994  ] =    292;
		rom[ 995  ] =    -63;
		rom[ 996  ] =    -10;
		rom[ 997  ] =    150;
		rom[ 998  ] =     39;
		rom[ 999  ] =     43;
		rom[ 1000 ] =    -38;
		rom[ 1001 ] =   -102;
		rom[ 1002 ] =     71;
		rom[ 1003 ] =      0;
		rom[ 1004 ] =    105;
		rom[ 1005 ] =   -365;
		rom[ 1006 ] =    -64;
		rom[ 1007 ] =     11;
		rom[ 1008 ] =   -240;
		rom[ 1009 ] =    -69;
		rom[ 1010 ] =   -264;
		rom[ 1011 ] =    161;
		rom[ 1012 ] =     41;
		rom[ 1013 ] =    -64;
		rom[ 1014 ] =    -74;
		rom[ 1015 ] =     -2;
		rom[ 1016 ] =     28;
		rom[ 1017 ] =    -49;
		rom[ 1018 ] =     79;
		rom[ 1019 ] =     -1;
		rom[ 1020 ] =   -117;
		rom[ 1021 ] =     -3;
		rom[ 1022 ] =    -19;
		rom[ 1023 ] =    -68;
		rom[ 1024 ] =     46;
		rom[ 1025 ] =    -48;
		rom[ 1026 ] =    -37;
		rom[ 1027 ] =   -134;
		rom[ 1028 ] =    -98;
		rom[ 1029 ] =     -1;
		rom[ 1030 ] =   -148;
		rom[ 1031 ] =      5;
		rom[ 1032 ] =   -166;
		rom[ 1033 ] =    -86;
		rom[ 1034 ] =     38;
		rom[ 1035 ] =    -64;
		rom[ 1036 ] =    -28;
		rom[ 1037 ] =   -249;
		rom[ 1038 ] =     97;
		rom[ 1039 ] =   -266;
		rom[ 1040 ] =  -1410;
		rom[ 1041 ] =    244;
		rom[ 1042 ] =      2;
		rom[ 1043 ] =     57;
		rom[ 1044 ] =     42;
		rom[ 1045 ] =   -221;
		rom[ 1046 ] =   -721;
		rom[ 1047 ] =   -331;
		rom[ 1048 ] =   -208;
		rom[ 1049 ] =    168;
		rom[ 1050 ] =      1;
		rom[ 1051 ] =     78;
		rom[ 1052 ] =     65;
		rom[ 1053 ] =   -367;
		rom[ 1054 ] =    -43;
		rom[ 1055 ] =   -166;
		rom[ 1056 ] =    -13;
		rom[ 1057 ] =   -235;
		rom[ 1058 ] =    137;
		rom[ 1059 ] =   -139;
		rom[ 1060 ] =     39;
		rom[ 1061 ] =    -62;
		rom[ 1062 ] =   -130;
		rom[ 1063 ] =    -55;
		rom[ 1064 ] =     29;
		rom[ 1065 ] =     -3;
		rom[ 1066 ] =    311;
		rom[ 1067 ] =    -64;
		rom[ 1068 ] =     57;
		rom[ 1069 ] =     64;
		rom[ 1070 ] =    -83;
		rom[ 1071 ] =    -14;
		rom[ 1072 ] =      0;
		rom[ 1073 ] =    -78;
		rom[ 1074 ] =    -62;
		rom[ 1075 ] =    120;
		rom[ 1076 ] =     98;
		rom[ 1077 ] =    -12;
		rom[ 1078 ] =     54;
		rom[ 1079 ] =    -43;
		rom[ 1080 ] =     29;
		rom[ 1081 ] =    -11;
		rom[ 1082 ] =   -103;
		rom[ 1083 ] =    -84;
		rom[ 1084 ] =   -185;
		rom[ 1085 ] =    -40;
		rom[ 1086 ] =     49;
		rom[ 1087 ] =    210;
		rom[ 1088 ] =   -110;
		rom[ 1089 ] =     -7;
		rom[ 1090 ] =     28;
		rom[ 1091 ] =    557;
		rom[ 1092 ] =    -12;
		rom[ 1093 ] =    -83;
		rom[ 1094 ] =    294;
		rom[ 1095 ] =    -99;
		rom[ 1096 ] =   -429;
		rom[ 1097 ] =   -249;
		rom[ 1098 ] =     53;
		rom[ 1099 ] =    -42;
		rom[ 1100 ] =     60;
		rom[ 1101 ] =   -237;
		rom[ 1102 ] =   -188;
		rom[ 1103 ] =     36;
		rom[ 1104 ] =      2;
		rom[ 1105 ] =   -304;
		rom[ 1106 ] =    622;
		rom[ 1107 ] =    183;
		rom[ 1108 ] =     40;
		rom[ 1109 ] =   -208;
		rom[ 1110 ] =    238;
		rom[ 1111 ] =   -144;
		rom[ 1112 ] =   -202;
		rom[ 1113 ] =   -362;
		rom[ 1114 ] =     97;
		rom[ 1115 ] =   -104;
		rom[ 1116 ] =    -61;
		rom[ 1117 ] =   -223;
		rom[ 1118 ] =     39;
		rom[ 1119 ] =   -293;
		rom[ 1120 ] =     39;
		rom[ 1121 ] =     10;
		rom[ 1122 ] =    111;
		rom[ 1123 ] =    111;
		rom[ 1124 ] =    -24;
		rom[ 1125 ] =    -97;
		rom[ 1126 ] =    228;
		rom[ 1127 ] =    220;
		rom[ 1128 ] =    153;
		rom[ 1129 ] =   -406;
		rom[ 1130 ] =     43;
		rom[ 1131 ] =    130;
		rom[ 1132 ] =   -110;
		rom[ 1133 ] =    -80;
		rom[ 1134 ] =    270;
		rom[ 1135 ] =   -183;
		rom[ 1136 ] =     63;
		rom[ 1137 ] =   -176;
		rom[ 1138 ] =   -151;
		rom[ 1139 ] =     11;
		rom[ 1140 ] =   -157;
		rom[ 1141 ] =    -78;
		rom[ 1142 ] =   -351;
		rom[ 1143 ] =   -143;
		rom[ 1144 ] =      1;
		rom[ 1145 ] =    400;
		rom[ 1146 ] =   -404;
		rom[ 1147 ] =   -397;
		rom[ 1148 ] =     44;
		rom[ 1149 ] =   -334;
		rom[ 1150 ] =   -353;
		rom[ 1151 ] =   -181;
		rom[ 1152 ] =    -10;
		rom[ 1153 ] =    147;
		rom[ 1154 ] =   -126;
		rom[ 1155 ] =   -125;
		rom[ 1156 ] =   -154;
		rom[ 1157 ] =     60;
		rom[ 1158 ] =    -20;
		rom[ 1159 ] =   -308;
		rom[ 1160 ] =     59;
		rom[ 1161 ] =   -207;
		rom[ 1162 ] =    157;
		rom[ 1163 ] =    -75;
		rom[ 1164 ] =   -156;
		rom[ 1165 ] =   -136;
		rom[ 1166 ] =   -329;
		rom[ 1167 ] =    -43;
		rom[ 1168 ] =    -28;
		rom[ 1169 ] =    261;
		rom[ 1170 ] =   -200;
		rom[ 1171 ] =   -225;
		rom[ 1172 ] =     29;
		rom[ 1173 ] =   -207;
		rom[ 1174 ] =    -18;
		rom[ 1175 ] =   -329;
		rom[ 1176 ] =    121;
		rom[ 1177 ] =    -15;
		rom[ 1178 ] =     44;
		rom[ 1179 ] =    -51;
		rom[ 1180 ] =    -17;
		rom[ 1181 ] =   -326;
		rom[ 1182 ] =     31;
		rom[ 1183 ] =      3;
		rom[ 1184 ] =    158;
		rom[ 1185 ] =    -92;
		rom[ 1186 ] =    134;
		rom[ 1187 ] =    -43;
		rom[ 1188 ] =   -304;
		rom[ 1189 ] =    214;
		rom[ 1190 ] =     90;
		rom[ 1191 ] =   -225;
		rom[ 1192 ] =    -36;
		rom[ 1193 ] =    -74;
		rom[ 1194 ] =     -8;
		rom[ 1195 ] =    177;
		rom[ 1196 ] =   -165;
		rom[ 1197 ] =     -7;
		rom[ 1198 ] =     -2;
		rom[ 1199 ] =    217;
		rom[ 1200 ] =   -531;
		rom[ 1201 ] =   -219;
		rom[ 1202 ] =     98;
		rom[ 1203 ] =   -441;
		rom[ 1204 ] =    140;
		rom[ 1205 ] =     -9;
		rom[ 1206 ] =    149;
		rom[ 1207 ] =     -3;
		rom[ 1208 ] =     38;
		rom[ 1209 ] =    132;
		rom[ 1210 ] =     -5;
		rom[ 1211 ] =   -220;
		rom[ 1212 ] =   -116;
		rom[ 1213 ] =     33;
		rom[ 1214 ] =     33;
		rom[ 1215 ] =    -64;
		rom[ 1216 ] =      5;
		rom[ 1217 ] =   -100;
		rom[ 1218 ] =     21;
		rom[ 1219 ] =    -46;
		rom[ 1220 ] =   -158;
		rom[ 1221 ] =    -12;
		rom[ 1222 ] =     45;
		rom[ 1223 ] =   -215;
		rom[ 1224 ] =    -48;
		rom[ 1225 ] =   -203;
		rom[ 1226 ] =    -60;
		rom[ 1227 ] =    -14;
		rom[ 1228 ] =     67;
		rom[ 1229 ] =   -171;
		rom[ 1230 ] =    172;
		rom[ 1231 ] =     77;
		rom[ 1232 ] =     37;
		rom[ 1233 ] =    -47;
		rom[ 1234 ] =     48;
		rom[ 1235 ] =    115;
		rom[ 1236 ] =     34;
		rom[ 1237 ] =    -53;
		rom[ 1238 ] =     82;
		rom[ 1239 ] =    -51;
		rom[ 1240 ] =     40;
		rom[ 1241 ] =   -160;
		rom[ 1242 ] =     42;
		rom[ 1243 ] =    -64;
		rom[ 1244 ] =     39;
		rom[ 1245 ] =    145;
		rom[ 1246 ] =    146;
		rom[ 1247 ] =    -98;
		rom[ 1248 ] =     56;
		rom[ 1249 ] =    -73;
		rom[ 1250 ] =   -166;
		rom[ 1251 ] =    -74;
		rom[ 1252 ] =    116;
		rom[ 1253 ] =   -131;
		rom[ 1254 ] =      4;
		rom[ 1255 ] =    100;
		rom[ 1256 ] =    304;
		rom[ 1257 ] =   -174;
		rom[ 1258 ] =   -217;
		rom[ 1259 ] =   -282;
		rom[ 1260 ] =    -50;
		rom[ 1261 ] =   -104;
		rom[ 1262 ] =    -75;
		rom[ 1263 ] =   -334;
		rom[ 1264 ] =     60;
		rom[ 1265 ] =     74;
		rom[ 1266 ] =   -620;
		rom[ 1267 ] =    225;
		rom[ 1268 ] =    205;
		rom[ 1269 ] =     37;
		rom[ 1270 ] =   -208;
		rom[ 1271 ] =   -181;
		rom[ 1272 ] =   -186;
		rom[ 1273 ] =     43;
		rom[ 1274 ] =    708;
		rom[ 1275 ] =     29;
		rom[ 1276 ] =     -1;
		rom[ 1277 ] =     59;
		rom[ 1278 ] =    -79;
		rom[ 1279 ] =    -12;
		rom[ 1280 ] =   -297;
		rom[ 1281 ] =    -69;
		rom[ 1282 ] =   -138;
		rom[ 1283 ] =     46;
		rom[ 1284 ] =    160;
		rom[ 1285 ] =     61;
		rom[ 1286 ] =   -240;
		rom[ 1287 ] =    -19;
		rom[ 1288 ] =     10;
		rom[ 1289 ] =     43;
		rom[ 1290 ] =     -8;
		rom[ 1291 ] =     24;
		rom[ 1292 ] =   -101;
		rom[ 1293 ] =    -58;
		rom[ 1294 ] =    -70;
		rom[ 1295 ] =    -27;
		rom[ 1296 ] =    -12;
		rom[ 1297 ] =     38;
		rom[ 1298 ] =     -5;
		rom[ 1299 ] =   -205;
		rom[ 1300 ] =    -53;
		rom[ 1301 ] =     51;
		rom[ 1302 ] =    -46;
		rom[ 1303 ] =    127;
		rom[ 1304 ] =    299;
		rom[ 1305 ] =    -16;
		rom[ 1306 ] =    -59;
		rom[ 1307 ] =   -210;
		rom[ 1308 ] =    155;
		rom[ 1309 ] =    -10;
		rom[ 1310 ] =   -294;
		rom[ 1311 ] =     -2;
		rom[ 1312 ] =     96;
		rom[ 1313 ] =    -25;
		rom[ 1314 ] =    171;
		rom[ 1315 ] =     40;
		rom[ 1316 ] =     97;
		rom[ 1317 ] =     38;
		rom[ 1318 ] =   -174;
		rom[ 1319 ] =     65;
		rom[ 1320 ] =     -7;
		rom[ 1321 ] =    -90;
		rom[ 1322 ] =     -9;
		rom[ 1323 ] =     -6;
		rom[ 1324 ] =     27;
		rom[ 1325 ] =    119;
		rom[ 1326 ] =    -72;
		rom[ 1327 ] =     -5;
		rom[ 1328 ] =    -83;
		rom[ 1329 ] =   -313;
		rom[ 1330 ] =     -4;
		rom[ 1331 ] =    167;
		rom[ 1332 ] =   -133;
		rom[ 1333 ] =   -200;
		rom[ 1334 ] =      0;
		rom[ 1335 ] =    -13;
		rom[ 1336 ] =      4;
		rom[ 1337 ] =   -159;
		rom[ 1338 ] =     45;
		rom[ 1339 ] =     11;
		rom[ 1340 ] =    116;
		rom[ 1341 ] =     85;
		rom[ 1342 ] =   -598;
		rom[ 1343 ] =   -169;
		rom[ 1344 ] =    117;
		rom[ 1345 ] =    -68;
		rom[ 1346 ] =    -47;
		rom[ 1347 ] =     -6;
		rom[ 1348 ] =     -8;
		rom[ 1349 ] =      1;
		rom[ 1350 ] =    108;
		rom[ 1351 ] =     -5;
		rom[ 1352 ] =     -8;
		rom[ 1353 ] =     28;
		rom[ 1354 ] =     74;
		rom[ 1355 ] =     30;
		rom[ 1356 ] =     37;
		rom[ 1357 ] =   -137;
		rom[ 1358 ] =    -15;
		rom[ 1359 ] =   -115;
		rom[ 1360 ] =    310;
		rom[ 1361 ] =   -590;
		rom[ 1362 ] =   -183;
		rom[ 1363 ] =     18;
		rom[ 1364 ] =   -313;
		rom[ 1365 ] =     34;
		rom[ 1366 ] =     -7;
		rom[ 1367 ] =     34;
		rom[ 1368 ] =    -37;
		rom[ 1369 ] =     49;
		rom[ 1370 ] =    -95;
		rom[ 1371 ] =    207;
		rom[ 1372 ] =    214;
		rom[ 1373 ] =   -242;
		rom[ 1374 ] =     11;
		rom[ 1375 ] =   -497;
		rom[ 1376 ] =    -54;
		rom[ 1377 ] =    153;
		rom[ 1378 ] =    -56;
		rom[ 1379 ] =    161;
		rom[ 1380 ] =    -59;
		rom[ 1381 ] =     46;
		rom[ 1382 ] =   -178;
		rom[ 1383 ] =     88;
		rom[ 1384 ] =   -224;
		rom[ 1385 ] =     60;
		rom[ 1386 ] =    -15;
		rom[ 1387 ] =    -50;
		rom[ 1388 ] =    247;
		rom[ 1389 ] =    -15;
		rom[ 1390 ] =   -116;
		rom[ 1391 ] =     29;
		rom[ 1392 ] =    463;
		rom[ 1393 ] =     59;
		rom[ 1394 ] =    126;
		rom[ 1395 ] =    155;
		rom[ 1396 ] =    102;
		rom[ 1397 ] =   -217;
		rom[ 1398 ] =   -202;
		rom[ 1399 ] =   -172;
		rom[ 1400 ] =      9;
		rom[ 1401 ] =     35;
		rom[ 1402 ] =    -35;
		rom[ 1403 ] =     35;
		rom[ 1404 ] =    -51;
		rom[ 1405 ] =   -119;
		rom[ 1406 ] =   -241;
		rom[ 1407 ] =     83;
		rom[ 1408 ] =     70;
		rom[ 1409 ] =     60;
		rom[ 1410 ] =   -147;
		rom[ 1411 ] =   -156;
		rom[ 1412 ] =   -144;
		rom[ 1413 ] =   -205;
		rom[ 1414 ] =   -207;
		rom[ 1415 ] =     35;
		rom[ 1416 ] =    -42;
		rom[ 1417 ] =    369;
		rom[ 1418 ] =     34;
		rom[ 1419 ] =    -86;
		rom[ 1420 ] =    -29;
		rom[ 1421 ] =   -254;
		rom[ 1422 ] =   -123;
		rom[ 1423 ] =      9;
		rom[ 1424 ] =   -278;
		rom[ 1425 ] =    244;
		rom[ 1426 ] =   -265;
		rom[ 1427 ] =    230;
		rom[ 1428 ] =   -259;
		rom[ 1429 ] =    157;
		rom[ 1430 ] =    -21;
		rom[ 1431 ] =     16;
		rom[ 1432 ] =   -239;
		rom[ 1433 ] =   -215;
		rom[ 1434 ] =    155;
		rom[ 1435 ] =     -7;
		rom[ 1436 ] =     33;
		rom[ 1437 ] =   -289;
		rom[ 1438 ] =    194;
		rom[ 1439 ] =     76;
		rom[ 1440 ] =      5;
		rom[ 1441 ] =   -218;
		rom[ 1442 ] =    -15;
		rom[ 1443 ] =     91;
		rom[ 1444 ] =      0;
		rom[ 1445 ] =     -8;
		rom[ 1446 ] =    151;
		rom[ 1447 ] =    152;
		rom[ 1448 ] =   -300;
		rom[ 1449 ] =     -4;
		rom[ 1450 ] =     41;
		rom[ 1451 ] =    -57;
		rom[ 1452 ] =     70;
		rom[ 1453 ] =   -194;
		rom[ 1454 ] =    -58;
		rom[ 1455 ] =     49;
		rom[ 1456 ] =     42;
		rom[ 1457 ] =    328;
		rom[ 1458 ] =   -138;
		rom[ 1459 ] =    162;
		rom[ 1460 ] =   -127;
		rom[ 1461 ] =   -303;
		rom[ 1462 ] =      5;
		rom[ 1463 ] =      7;
		rom[ 1464 ] =    -53;
		rom[ 1465 ] =      0;
		rom[ 1466 ] =    -56;
		rom[ 1467 ] =     -2;
		rom[ 1468 ] =    114;
		rom[ 1469 ] =    -52;
		rom[ 1470 ] =   -196;
		rom[ 1471 ] =   -361;
		rom[ 1472 ] =     49;
		rom[ 1473 ] =    215;
		rom[ 1474 ] =     32;
		rom[ 1475 ] =   -119;
		rom[ 1476 ] =    132;
		rom[ 1477 ] =     -7;
		rom[ 1478 ] =     62;
		rom[ 1479 ] =    250;
		rom[ 1480 ] =     51;
		rom[ 1481 ] =    -65;
		rom[ 1482 ] =     43;
		rom[ 1483 ] =   -219;
		rom[ 1484 ] =    143;
		rom[ 1485 ] =    -65;
		rom[ 1486 ] =      1;
		rom[ 1487 ] =   -154;
		rom[ 1488 ] =    107;
		rom[ 1489 ] =     58;
		rom[ 1490 ] =     23;
		rom[ 1491 ] =    -68;
		rom[ 1492 ] =   -185;
		rom[ 1493 ] =    -89;
		rom[ 1494 ] =     29;
		rom[ 1495 ] =     -2;
		rom[ 1496 ] =     52;
		rom[ 1497 ] =    148;
		rom[ 1498 ] =      4;
		rom[ 1499 ] =    -84;
		rom[ 1500 ] =    351;
		rom[ 1501 ] =      0;
		rom[ 1502 ] =     -3;
		rom[ 1503 ] =     96;
		rom[ 1504 ] =   -703;
		rom[ 1505 ] =    121;
		rom[ 1506 ] =   -148;
		rom[ 1507 ] =     -2;
		rom[ 1508 ] =     89;
		rom[ 1509 ] =    364;
		rom[ 1510 ] =     61;
		rom[ 1511 ] =     -2;
		rom[ 1512 ] =     -4;
		rom[ 1513 ] =   -231;
		rom[ 1514 ] =    -54;
		rom[ 1515 ] =     50;
		rom[ 1516 ] =    -23;
		rom[ 1517 ] =   -141;
		rom[ 1518 ] =     47;
		rom[ 1519 ] =    496;
		rom[ 1520 ] =    -67;
		rom[ 1521 ] =   -140;
		rom[ 1522 ] =   -655;
		rom[ 1523 ] =    -63;
		rom[ 1524 ] =     41;
		rom[ 1525 ] =     56;
		rom[ 1526 ] =     79;
		rom[ 1527 ] =   -244;
		rom[ 1528 ] =     32;
		rom[ 1529 ] =    -15;
		rom[ 1530 ] =     10;
		rom[ 1531 ] =    -11;
		rom[ 1532 ] =     10;
		rom[ 1533 ] =      7;
		rom[ 1534 ] =    264;
		rom[ 1535 ] =    -17;
		rom[ 1536 ] =   -152;
		rom[ 1537 ] =    -16;
		rom[ 1538 ] =     14;
		rom[ 1539 ] =     -1;
		rom[ 1540 ] =     37;
		rom[ 1541 ] =    -45;
		rom[ 1542 ] =   -152;
		rom[ 1543 ] =   -276;
		rom[ 1544 ] =    199;
		rom[ 1545 ] =    -16;
		rom[ 1546 ] =     -4;
		rom[ 1547 ] =    -14;
		rom[ 1548 ] =     87;
		rom[ 1549 ] =    -67;
		rom[ 1550 ] =    -33;
		rom[ 1551 ] =      7;
		rom[ 1552 ] =      6;
		rom[ 1553 ] =    115;
		rom[ 1554 ] =    -50;
		rom[ 1555 ] =   -138;
		rom[ 1556 ] =     -3;
		rom[ 1557 ] =     17;
		rom[ 1558 ] =    174;
		rom[ 1559 ] =    -52;
		rom[ 1560 ] =    182;
		rom[ 1561 ] =    -94;
		rom[ 1562 ] =   -220;
		rom[ 1563 ] =    -69;
		rom[ 1564 ] =    -88;
		rom[ 1565 ] =    -81;
		rom[ 1566 ] =   -176;
		rom[ 1567 ] =    -53;
		rom[ 1568 ] =   -126;
		rom[ 1569 ] =    343;
		rom[ 1570 ] =     11;
		rom[ 1571 ] =   -182;
		rom[ 1572 ] =    257;
		rom[ 1573 ] =     -3;
		rom[ 1574 ] =   -209;
		rom[ 1575 ] =    138;
		rom[ 1576 ] =    -86;
		rom[ 1577 ] =   -306;
		rom[ 1578 ] =   -227;
		rom[ 1579 ] =     42;
		rom[ 1580 ] =    160;
		rom[ 1581 ] =    -72;
		rom[ 1582 ] =   -163;
		rom[ 1583 ] =   -196;
		rom[ 1584 ] =    116;
		rom[ 1585 ] =   -195;
		rom[ 1586 ] =     11;
		rom[ 1587 ] =    -12;
		rom[ 1588 ] =     -5;
		rom[ 1589 ] =   -245;
		rom[ 1590 ] =   -179;
		rom[ 1591 ] =    -72;
		rom[ 1592 ] =    -64;
		rom[ 1593 ] =   -178;
		rom[ 1594 ] =    117;
		rom[ 1595 ] =     46;
		rom[ 1596 ] =   -161;
		rom[ 1597 ] =   -263;
		rom[ 1598 ] =     88;
		rom[ 1599 ] =    -74;
		rom[ 1600 ] =   -113;
		rom[ 1601 ] =     45;
		rom[ 1602 ] =     -2;
		rom[ 1603 ] =    423;
		rom[ 1604 ] =     -1;
		rom[ 1605 ] =      0;
		rom[ 1606 ] =   -158;
		rom[ 1607 ] =    180;
		rom[ 1608 ] =    100;
		rom[ 1609 ] =     -6;
		rom[ 1610 ] =    120;
		rom[ 1611 ] =     82;
		rom[ 1612 ] =   -314;
		rom[ 1613 ] =     11;
		rom[ 1614 ] =    -42;
		rom[ 1615 ] =     86;
		rom[ 1616 ] =   -218;
		rom[ 1617 ] =     14;
		rom[ 1618 ] =    133;
		rom[ 1619 ] =    160;
		rom[ 1620 ] =   -157;
		rom[ 1621 ] =   -216;
		rom[ 1622 ] =    -16;
		rom[ 1623 ] =    -45;
		rom[ 1624 ] =     -7;
		rom[ 1625 ] =    -62;
		rom[ 1626 ] =    -60;
		rom[ 1627 ] =    100;
		rom[ 1628 ] =    -68;
		rom[ 1629 ] =     44;
		rom[ 1630 ] =   -277;
		rom[ 1631 ] =    184;
		rom[ 1632 ] =   -304;
		rom[ 1633 ] =    161;
		rom[ 1634 ] =    338;
		rom[ 1635 ] =    -86;
		rom[ 1636 ] =    -65;
		rom[ 1637 ] =     36;
		rom[ 1638 ] =   -298;
		rom[ 1639 ] =   -101;
		rom[ 1640 ] =    126;
		rom[ 1641 ] =    479;
		rom[ 1642 ] =   -227;
		rom[ 1643 ] =   -298;
		rom[ 1644 ] =   -171;
		rom[ 1645 ] =   -122;
		rom[ 1646 ] =     30;
		rom[ 1647 ] =    -19;
		rom[ 1648 ] =    -51;
		rom[ 1649 ] =    236;
		rom[ 1650 ] =    -68;
		rom[ 1651 ] =   -138;
		rom[ 1652 ] =      4;
		rom[ 1653 ] =     -3;
		rom[ 1654 ] =    -45;
		rom[ 1655 ] =     53;
		rom[ 1656 ] =      5;
		rom[ 1657 ] =     -4;
		rom[ 1658 ] =    -48;
		rom[ 1659 ] =    104;
		rom[ 1660 ] =    -52;
		rom[ 1661 ] =   -434;
		rom[ 1662 ] =     -7;
		rom[ 1663 ] =    -51;
		rom[ 1664 ] =   -115;
		rom[ 1665 ] =     60;
		rom[ 1666 ] =    -46;
		rom[ 1667 ] =    -70;
		rom[ 1668 ] =   -118;
		rom[ 1669 ] =    106;
		rom[ 1670 ] =     37;
		rom[ 1671 ] =    192;
		rom[ 1672 ] =    -48;
		rom[ 1673 ] =     90;
		rom[ 1674 ] =   -164;
		rom[ 1675 ] =      4;
		rom[ 1676 ] =    270;
		rom[ 1677 ] =     76;
		rom[ 1678 ] =    -55;
		rom[ 1679 ] =     61;
		rom[ 1680 ] =     -8;
		rom[ 1681 ] =     -1;
		rom[ 1682 ] =     19;
		rom[ 1683 ] =     20;
		rom[ 1684 ] =    -35;
		rom[ 1685 ] =   -476;
		rom[ 1686 ] =    -47;
		rom[ 1687 ] =     36;
		rom[ 1688 ] =    411;
		rom[ 1689 ] =   -207;
		rom[ 1690 ] =   -356;
		rom[ 1691 ] =      8;
		rom[ 1692 ] =   -141;
		rom[ 1693 ] =      5;
		rom[ 1694 ] =    113;
		rom[ 1695 ] =     46;
		rom[ 1696 ] =    -16;
		rom[ 1697 ] =     51;
		rom[ 1698 ] =    -81;
		rom[ 1699 ] =    222;
		rom[ 1700 ] =    163;
		rom[ 1701 ] =     44;
		rom[ 1702 ] =     61;
		rom[ 1703 ] =    138;
		rom[ 1704 ] =    612;
		rom[ 1705 ] =     40;
		rom[ 1706 ] =      0;
		rom[ 1707 ] =    -29;
		rom[ 1708 ] =   -269;
		rom[ 1709 ] =    -51;
		rom[ 1710 ] =    -54;
		rom[ 1711 ] =     28;
		rom[ 1712 ] =   -439;
		rom[ 1713 ] =    165;
		rom[ 1714 ] =     -2;
		rom[ 1715 ] =     50;
		rom[ 1716 ] =   -221;
		rom[ 1717 ] =     35;
		rom[ 1718 ] =     86;
		rom[ 1719 ] =   -640;
		rom[ 1720 ] =    129;
		rom[ 1721 ] =   -750;
		rom[ 1722 ] =   -153;
		rom[ 1723 ] =     86;
		rom[ 1724 ] =   -283;
		rom[ 1725 ] =    114;
		rom[ 1726 ] =   -266;
		rom[ 1727 ] =      8;
		rom[ 1728 ] =    135;
		rom[ 1729 ] =   -137;
		rom[ 1730 ] =   -128;
		rom[ 1731 ] =    -84;
		rom[ 1732 ] =    -81;
		rom[ 1733 ] =     27;
		rom[ 1734 ] =    -36;
		rom[ 1735 ] =    241;
		rom[ 1736 ] =   -139;
		rom[ 1737 ] =      3;
		rom[ 1738 ] =    -80;
		rom[ 1739 ] =     -1;
		rom[ 1740 ] =   -195;
		rom[ 1741 ] =     61;
		rom[ 1742 ] =    -24;
		rom[ 1743 ] =   -202;
		rom[ 1744 ] =    -26;
		rom[ 1745 ] =   -103;
		rom[ 1746 ] =     52;
		rom[ 1747 ] =      0;
		rom[ 1748 ] =     -1;
		rom[ 1749 ] =    -93;
		rom[ 1750 ] =   -365;
		rom[ 1751 ] =    -10;
		rom[ 1752 ] =     67;
		rom[ 1753 ] =   -214;
		rom[ 1754 ] =   -125;
		rom[ 1755 ] =    -48;
		rom[ 1756 ] =     59;
		rom[ 1757 ] =     -9;
		rom[ 1758 ] =   -456;
		rom[ 1759 ] =    -55;
		rom[ 1760 ] =    -45;
		rom[ 1761 ] =     -2;
		rom[ 1762 ] =     77;
		rom[ 1763 ] =   -243;
		rom[ 1764 ] =      8;
		rom[ 1765 ] =    250;
		rom[ 1766 ] =     -5;
		rom[ 1767 ] =    -14;
		rom[ 1768 ] =    167;
		rom[ 1769 ] =      6;
		rom[ 1770 ] =     -1;
		rom[ 1771 ] =     87;
		rom[ 1772 ] =     -1;
		rom[ 1773 ] =   -134;
		rom[ 1774 ] =   -149;
		rom[ 1775 ] =      5;
		rom[ 1776 ] =    -93;
		rom[ 1777 ] =      9;
		rom[ 1778 ] =    -37;
		rom[ 1779 ] =    -55;
		rom[ 1780 ] =   -277;
		rom[ 1781 ] =    -39;
		rom[ 1782 ] =     11;
		rom[ 1783 ] =   -396;
		rom[ 1784 ] =     42;
		rom[ 1785 ] =   -197;
		rom[ 1786 ] =     28;
		rom[ 1787 ] =    283;
		rom[ 1788 ] =     70;
		rom[ 1789 ] =   -206;
		rom[ 1790 ] =     36;
		rom[ 1791 ] =     50;
		rom[ 1792 ] =    -12;
		rom[ 1793 ] =    -42;
		rom[ 1794 ] =    -32;
		rom[ 1795 ] =     -8;
		rom[ 1796 ] =    -16;
		rom[ 1797 ] =    -93;
		rom[ 1798 ] =     30;
		rom[ 1799 ] =   -133;
		rom[ 1800 ] =    166;
		rom[ 1801 ] =     44;
		rom[ 1802 ] =    -50;
		rom[ 1803 ] =   -130;
		rom[ 1804 ] =    -17;
		rom[ 1805 ] =   -104;
		rom[ 1806 ] =    -54;
		rom[ 1807 ] =   -127;
		rom[ 1808 ] =    -52;
		rom[ 1809 ] =     46;
		rom[ 1810 ] =      3;
		rom[ 1811 ] =    -53;
		rom[ 1812 ] =     63;
		rom[ 1813 ] =   -488;
		rom[ 1814 ] =   -182;
		rom[ 1815 ] =    -43;
		rom[ 1816 ] =     48;
		rom[ 1817 ] =      1;
		rom[ 1818 ] =     43;
		rom[ 1819 ] =   -578;
		rom[ 1820 ] =    616;
		rom[ 1821 ] =    -69;
		rom[ 1822 ] =     80;
		rom[ 1823 ] =   -371;
		rom[ 1824 ] =     -4;
		rom[ 1825 ] =    -59;
		rom[ 1826 ] =     36;
		rom[ 1827 ] =    -56;
		rom[ 1828 ] =    -29;
		rom[ 1829 ] =      6;
		rom[ 1830 ] =     45;
		rom[ 1831 ] =    -37;
		rom[ 1832 ] =   -134;
		rom[ 1833 ] =    225;
		rom[ 1834 ] =   -123;
		rom[ 1835 ] =    -54;
		rom[ 1836 ] =    -18;
		rom[ 1837 ] =    -63;
		rom[ 1838 ] =      2;
		rom[ 1839 ] =    -45;
		rom[ 1840 ] =     33;
		rom[ 1841 ] =    -11;
		rom[ 1842 ] =     44;
		rom[ 1843 ] =   -289;
		rom[ 1844 ] =    -57;
		rom[ 1845 ] =    116;
		rom[ 1846 ] =    -38;
		rom[ 1847 ] =   -174;
		rom[ 1848 ] =    166;
		rom[ 1849 ] =    114;
		rom[ 1850 ] =    -22;
		rom[ 1851 ] =   -119;
		rom[ 1852 ] =     74;
		rom[ 1853 ] =   -309;
		rom[ 1854 ] =    -11;
		rom[ 1855 ] =    -68;
		rom[ 1856 ] =    -33;
		rom[ 1857 ] =    497;
		rom[ 1858 ] =     39;
		rom[ 1859 ] =   -182;
		rom[ 1860 ] =    235;
		rom[ 1861 ] =    -57;
		rom[ 1862 ] =   -185;
		rom[ 1863 ] =    319;
		rom[ 1864 ] =   -370;
		rom[ 1865 ] =   -200;
		rom[ 1866 ] =   -218;
		rom[ 1867 ] =    -38;
		rom[ 1868 ] =    140;
		rom[ 1869 ] =     93;
		rom[ 1870 ] =     -8;
		rom[ 1871 ] =   -157;
		rom[ 1872 ] =    -16;
		rom[ 1873 ] =    -87;
		rom[ 1874 ] =    -77;
		rom[ 1875 ] =     19;
		rom[ 1876 ] =   -249;
		rom[ 1877 ] =     47;
		rom[ 1878 ] =    -15;
		rom[ 1879 ] =     83;
		rom[ 1880 ] =    -75;
		rom[ 1881 ] =   -310;
		rom[ 1882 ] =     33;
		rom[ 1883 ] =   -169;
		rom[ 1884 ] =     42;
		rom[ 1885 ] =    -13;
		rom[ 1886 ] =     51;
		rom[ 1887 ] =   -201;
		rom[ 1888 ] =     73;
		rom[ 1889 ] =    442;
		rom[ 1890 ] =      4;
		rom[ 1891 ] =    -19;
		rom[ 1892 ] =     81;
		rom[ 1893 ] =    196;
		rom[ 1894 ] =     47;
		rom[ 1895 ] =    -60;
		rom[ 1896 ] =     44;
		rom[ 1897 ] =    -11;
		rom[ 1898 ] =    205;
		rom[ 1899 ] =   -209;
		rom[ 1900 ] =     38;
		rom[ 1901 ] =   -186;
		rom[ 1902 ] =    145;
		rom[ 1903 ] =     10;
		rom[ 1904 ] =   -507;
		rom[ 1905 ] =    128;
		rom[ 1906 ] =    102;
		rom[ 1907 ] =   -196;
		rom[ 1908 ] =    221;
		rom[ 1909 ] =   -143;
		rom[ 1910 ] =     10;
		rom[ 1911 ] =    -49;
		rom[ 1912 ] =     47;
		rom[ 1913 ] =    -12;
		rom[ 1914 ] =    362;
		rom[ 1915 ] =    337;
		rom[ 1916 ] =     12;
		rom[ 1917 ] =    -53;
		rom[ 1918 ] =   -319;
		rom[ 1919 ] =     66;
		rom[ 1920 ] =     58;
		rom[ 1921 ] =   -220;
		rom[ 1922 ] =     80;
		rom[ 1923 ] =     64;
		rom[ 1924 ] =     68;
		rom[ 1925 ] =   -138;
		rom[ 1926 ] =    183;
		rom[ 1927 ] =   -149;
		rom[ 1928 ] =   -190;
		rom[ 1929 ] =     45;
		rom[ 1930 ] =   -275;
		rom[ 1931 ] =      6;
		rom[ 1932 ] =   -115;
		rom[ 1933 ] =    -69;
		rom[ 1934 ] =   -125;
		rom[ 1935 ] =    106;
		rom[ 1936 ] =     41;
		rom[ 1937 ] =   -282;
		rom[ 1938 ] =    166;
		rom[ 1939 ] =    107;
		rom[ 1940 ] =     90;
		rom[ 1941 ] =    -74;
		rom[ 1942 ] =   -338;
		rom[ 1943 ] =   -224;
		rom[ 1944 ] =     66;
		rom[ 1945 ] =   -253;
		rom[ 1946 ] =    162;
		rom[ 1947 ] =      6;
		rom[ 1948 ] =   -144;
		rom[ 1949 ] =      0;
		rom[ 1950 ] =    -24;
		rom[ 1951 ] =   -167;
		rom[ 1952 ] =   -119;
		rom[ 1953 ] =   -271;
		rom[ 1954 ] =    129;
		rom[ 1955 ] =    -78;
		rom[ 1956 ] =   -285;
		rom[ 1957 ] =   -222;
		rom[ 1958 ] =    168;
		rom[ 1959 ] =    -58;
		rom[ 1960 ] =     46;
		rom[ 1961 ] =    -84;
		rom[ 1962 ] =    -30;
		rom[ 1963 ] =     98;
		rom[ 1964 ] =   -228;
		rom[ 1965 ] =    137;
		rom[ 1966 ] =    -14;
		rom[ 1967 ] =   -390;
		rom[ 1968 ] =     19;
		rom[ 1969 ] =    -50;
		rom[ 1970 ] =   -163;
		rom[ 1971 ] =     21;
		rom[ 1972 ] =   -110;
		rom[ 1973 ] =    102;
		rom[ 1974 ] =    135;
		rom[ 1975 ] =    -99;
		rom[ 1976 ] =    224;
		rom[ 1977 ] =   -298;
		rom[ 1978 ] =    279;
		rom[ 1979 ] =     35;
		rom[ 1980 ] =     34;
		rom[ 1981 ] =     -3;
		rom[ 1982 ] =     45;
		rom[ 1983 ] =   -135;
		rom[ 1984 ] =    -28;
		rom[ 1985 ] =    100;
		rom[ 1986 ] =    -65;
		rom[ 1987 ] =     -6;
		rom[ 1988 ] =    202;
		rom[ 1989 ] =   -122;
		rom[ 1990 ] =    -44;
		rom[ 1991 ] =      0;
		rom[ 1992 ] =      4;
		rom[ 1993 ] =     51;
		rom[ 1994 ] =     47;
		rom[ 1995 ] =    -15;
		rom[ 1996 ] =    -83;
		rom[ 1997 ] =   -159;
		rom[ 1998 ] =     -8;
		rom[ 1999 ] =     50;
		rom[ 2000 ] =     52;
		rom[ 2001 ] =   -145;
		rom[ 2002 ] =    191;
		rom[ 2003 ] =    217;
		rom[ 2004 ] =     42;
		rom[ 2005 ] =   -340;
		rom[ 2006 ] =    -15;
		rom[ 2007 ] =    195;
		rom[ 2008 ] =     57;
		rom[ 2009 ] =   -407;
		rom[ 2010 ] =     30;
		rom[ 2011 ] =   -335;
		rom[ 2012 ] =      0;
		rom[ 2013 ] =    167;
		rom[ 2014 ] =     18;
		rom[ 2015 ] =   -172;
		rom[ 2016 ] =     85;
		rom[ 2017 ] =    116;
		rom[ 2018 ] =    -11;
		rom[ 2019 ] =     68;
		rom[ 2020 ] =   -212;
		rom[ 2021 ] =   -172;
		rom[ 2022 ] =    -18;
		rom[ 2023 ] =      7;
		rom[ 2024 ] =     34;
		rom[ 2025 ] =   -152;
		rom[ 2026 ] =    103;
		rom[ 2027 ] =   -278;
		rom[ 2028 ] =     74;
		rom[ 2029 ] =    167;
		rom[ 2030 ] =   -501;
		rom[ 2031 ] =    -58;
		rom[ 2032 ] =     40;
		rom[ 2033 ] =    -99;
		rom[ 2034 ] =    439;
		rom[ 2035 ] =    -97;
		rom[ 2036 ] =   -791;
		rom[ 2037 ] =    -35;
		rom[ 2038 ] =    -16;
		rom[ 2039 ] =   -144;
		rom[ 2040 ] =     64;
		rom[ 2041 ] =   -670;
		rom[ 2042 ] =     15;
		rom[ 2043 ] =    239;
		rom[ 2044 ] =     35;
		rom[ 2045 ] =     -3;
		rom[ 2046 ] =     15;
		rom[ 2047 ] =    182;
		rom[ 2048 ] =     37;
		rom[ 2049 ] =    -95;
		rom[ 2050 ] =    -60;
		rom[ 2051 ] =     -7;
		rom[ 2052 ] =     47;
		rom[ 2053 ] =    -39;
		rom[ 2054 ] =     38;
		rom[ 2055 ] =    -42;
		rom[ 2056 ] =    -18;
		rom[ 2057 ] =     -5;
		rom[ 2058 ] =    -46;
		rom[ 2059 ] =   -116;
		rom[ 2060 ] =     68;
		rom[ 2061 ] =    -39;
		rom[ 2062 ] =     17;
		rom[ 2063 ] =     70;
		rom[ 2064 ] =   -787;
		rom[ 2065 ] =   -374;
		rom[ 2066 ] =    226;
		rom[ 2067 ] =     35;
		rom[ 2068 ] =   -263;
		rom[ 2069 ] =     19;
		rom[ 2070 ] =     30;
		rom[ 2071 ] =    172;
		rom[ 2072 ] =     54;
		rom[ 2073 ] =    114;
		rom[ 2074 ] =      9;
		rom[ 2075 ] =    -50;
		rom[ 2076 ] =     34;
		rom[ 2077 ] =    215;
		rom[ 2078 ] =     44;
		rom[ 2079 ] =    -45;
		rom[ 2080 ] =    -36;
		rom[ 2081 ] =    267;
		rom[ 2082 ] =     28;
		rom[ 2083 ] =   -201;
		rom[ 2084 ] =   -155;
		rom[ 2085 ] =     -3;
		rom[ 2086 ] =   -523;
		rom[ 2087 ] =   -107;
		rom[ 2088 ] =      6;
		rom[ 2089 ] =    -44;
		rom[ 2090 ] =    -56;
		rom[ 2091 ] =    -17;
		rom[ 2092 ] =    330;
		rom[ 2093 ] =   -297;
		rom[ 2094 ] =     17;
		rom[ 2095 ] =    -45;
		rom[ 2096 ] =     56;
		rom[ 2097 ] =    158;
		rom[ 2098 ] =   -118;
		rom[ 2099 ] =    -32;
		rom[ 2100 ] =    -77;
		rom[ 2101 ] =    -57;
		rom[ 2102 ] =     64;
		rom[ 2103 ] =     74;
		rom[ 2104 ] =     49;
		rom[ 2105 ] =   -193;
		rom[ 2106 ] =     21;
		rom[ 2107 ] =    -68;
		rom[ 2108 ] =     34;
		rom[ 2109 ] =   -103;
		rom[ 2110 ] =     41;
		rom[ 2111 ] =     79;
		rom[ 2112 ] =    -68;
		rom[ 2113 ] =     39;
		rom[ 2114 ] =    293;
		rom[ 2115 ] =   -182;
		rom[ 2116 ] =    106;
		rom[ 2117 ] =   -341;
		rom[ 2118 ] =     36;
		rom[ 2119 ] =    -12;
		rom[ 2120 ] =    163;
		rom[ 2121 ] =    -55;
		rom[ 2122 ] =   -206;
		rom[ 2123 ] =    -81;
		rom[ 2124 ] =   -164;
		rom[ 2125 ] =   -117;
		rom[ 2126 ] =    117;
		rom[ 2127 ] =     93;
		rom[ 2128 ] =      6;
		rom[ 2129 ] =     44;
		rom[ 2130 ] =   -246;
		rom[ 2131 ] =   -181;
		rom[ 2132 ] =     18;
		rom[ 2133 ] =   -191;
		rom[ 2134 ] =    174;
		rom[ 2135 ] =    -32;
		rom[ 2136 ] =     18;
		rom[ 2137 ] =    244;
		rom[ 2138 ] =    -72;
		rom[ 2139 ] =     98;
		rom[ 2140 ] =      0;
		rom[ 2141 ] =    217;
		rom[ 2142 ] =   -236;
		rom[ 2143 ] =   -139;
		rom[ 2144 ] =     -1;
		rom[ 2145 ] =    184;
		rom[ 2146 ] =     49;
		rom[ 2147 ] =     29;
		rom[ 2148 ] =    -13;
		rom[ 2149 ] =    -27;
		rom[ 2150 ] =    -46;
		rom[ 2151 ] =     42;
		rom[ 2152 ] =     52;
		rom[ 2153 ] =    239;
		rom[ 2154 ] =      0;
		rom[ 2155 ] =      0;
		rom[ 2156 ] =    185;
		rom[ 2157 ] =    256;
		rom[ 2158 ] =    -11;
		rom[ 2159 ] =      3;
		rom[ 2160 ] =   -241;
		rom[ 2161 ] =   -111;
		rom[ 2162 ] =    -45;
		rom[ 2163 ] =    148;
		rom[ 2164 ] =     -5;
		rom[ 2165 ] =    -36;
		rom[ 2166 ] =    249;
		rom[ 2167 ] =    -21;
		rom[ 2168 ] =   -529;
		rom[ 2169 ] =    112;
		rom[ 2170 ] =     73;
		rom[ 2171 ] =   -146;
		rom[ 2172 ] =     88;
		rom[ 2173 ] =    143;
		rom[ 2174 ] =    -37;
		rom[ 2175 ] =     61;
		rom[ 2176 ] =    110;
		rom[ 2177 ] =      5;
		rom[ 2178 ] =     46;
		rom[ 2179 ] =     38;
		rom[ 2180 ] =    -50;
		rom[ 2181 ] =      0;
		rom[ 2182 ] =    323;
		rom[ 2183 ] =    166;
		rom[ 2184 ] =   -264;
		rom[ 2185 ] =   -122;
		rom[ 2186 ] =    -53;
		rom[ 2187 ] =    132;
		rom[ 2188 ] =    -54;
		rom[ 2189 ] =     46;
		rom[ 2190 ] =    -37;
		rom[ 2191 ] =    -72;
		rom[ 2192 ] =   -114;
		rom[ 2193 ] =     10;
		rom[ 2194 ] =    101;
		rom[ 2195 ] =    563;
		rom[ 2196 ] =    -71;
		rom[ 2197 ] =     87;
		rom[ 2198 ] =     73;
		rom[ 2199 ] =    163;
		rom[ 2200 ] =     20;
		rom[ 2201 ] =   -114;
		rom[ 2202 ] =   -251;
		rom[ 2203 ] =     58;
		rom[ 2204 ] =    214;
		rom[ 2205 ] =     29;
		rom[ 2206 ] =     -9;
		rom[ 2207 ] =   -346;
		rom[ 2208 ] =    -45;
		rom[ 2209 ] =     32;
		rom[ 2210 ] =    205;
		rom[ 2211 ] =     41;
		rom[ 2212 ] =     39;
		rom[ 2213 ] =   -471;
		rom[ 2214 ] =   -206;
		rom[ 2215 ] =    -35;
		rom[ 2216 ] =     -6;
		rom[ 2217 ] =   -188;
		rom[ 2218 ] =   -116;
		rom[ 2219 ] =     53;
		rom[ 2220 ] =    102;
		rom[ 2221 ] =     -5;
		rom[ 2222 ] =   -127;
		rom[ 2223 ] =     45;
		rom[ 2224 ] =     11;
		rom[ 2225 ] =     44;
		rom[ 2226 ] =   -118;
		rom[ 2227 ] =     13;
		rom[ 2228 ] =     38;
		rom[ 2229 ] =     35;
		rom[ 2230 ] =    -73;
		rom[ 2231 ] =    -77;
		rom[ 2232 ] =   -251;
		rom[ 2233 ] =     12;
		rom[ 2234 ] =     60;
		rom[ 2235 ] =    120;
		rom[ 2236 ] =    -53;
		rom[ 2237 ] =     42;
		rom[ 2238 ] =   -144;
		rom[ 2239 ] =   -911;
		rom[ 2240 ] =     -9;
		rom[ 2241 ] =   -144;
		rom[ 2242 ] =     -7;
		rom[ 2243 ] =   -136;
		rom[ 2244 ] =    -56;
		rom[ 2245 ] =     36;
		rom[ 2246 ] =    -88;
		rom[ 2247 ] =    245;
		rom[ 2248 ] =    445;
		rom[ 2249 ] =    355;
		rom[ 2250 ] =     13;
		rom[ 2251 ] =    -23;
		rom[ 2252 ] =      9;
		rom[ 2253 ] =    243;
		rom[ 2254 ] =    -34;
		rom[ 2255 ] =     58;
		rom[ 2256 ] =    -56;
		rom[ 2257 ] =    329;
		rom[ 2258 ] =  -1012;
		rom[ 2259 ] =     96;
		rom[ 2260 ] =     -6;
		rom[ 2261 ] =     43;
		rom[ 2262 ] =   -239;
		rom[ 2263 ] =     33;
		rom[ 2264 ] =   -292;
		rom[ 2265 ] =    126;
		rom[ 2266 ] =    -79;
		rom[ 2267 ] =    -97;
		rom[ 2268 ] =    -47;
		rom[ 2269 ] =   -151;
		rom[ 2270 ] =    -39;
		rom[ 2271 ] =     82;
		rom[ 2272 ] =    -40;
		rom[ 2273 ] =    193;
		rom[ 2274 ] =   -226;
		rom[ 2275 ] =     61;
		rom[ 2276 ] =   -479;
		rom[ 2277 ] =     33;
		rom[ 2278 ] =     -6;
		rom[ 2279 ] =    119;
		rom[ 2280 ] =    102;
		rom[ 2281 ] =   -400;
		rom[ 2282 ] =   -492;
		rom[ 2283 ] =     34;
		rom[ 2284 ] =    261;
		rom[ 2285 ] =    -24;
		rom[ 2286 ] =     28;
		rom[ 2287 ] =    154;
		rom[ 2288 ] =    -48;
		rom[ 2289 ] =     29;
		rom[ 2290 ] =    -71;
		rom[ 2291 ] =    185;
		rom[ 2292 ] =    -49;
		rom[ 2293 ] =     39;
		rom[ 2294 ] =    -14;
		rom[ 2295 ] =   -412;
		rom[ 2296 ] =    -15;
		rom[ 2297 ] =     41;
		rom[ 2298 ] =    -45;
		rom[ 2299 ] =   1190;
		rom[ 2300 ] =    -43;
		rom[ 2301 ] =    233;
		rom[ 2302 ] =     56;
		rom[ 2303 ] =   -230;
		rom[ 2304 ] =    -96;
		rom[ 2305 ] =    -97;
		rom[ 2306 ] =    -46;
		rom[ 2307 ] =    -57;
		rom[ 2308 ] =    181;
		rom[ 2309 ] =    122;
		rom[ 2310 ] =    -47;
		rom[ 2311 ] =     10;
		rom[ 2312 ] =    -59;
		rom[ 2313 ] =   -117;
		rom[ 2314 ] =     85;
		rom[ 2315 ] =    -42;
		rom[ 2316 ] =     57;
		rom[ 2317 ] =     38;
		rom[ 2318 ] =   -380;
		rom[ 2319 ] =    -49;
		rom[ 2320 ] =     34;
		rom[ 2321 ] =   -277;
		rom[ 2322 ] =   -151;
		rom[ 2323 ] =   -125;
		rom[ 2324 ] =    152;
		rom[ 2325 ] =   -302;
		rom[ 2326 ] =   -156;
		rom[ 2327 ] =   -292;
		rom[ 2328 ] =   -421;
		rom[ 2329 ] =    -79;
		rom[ 2330 ] =   -177;
		rom[ 2331 ] =   -183;
		rom[ 2332 ] =     57;
		rom[ 2333 ] =    264;
		rom[ 2334 ] =    115;
		rom[ 2335 ] =   -218;
		rom[ 2336 ] =    148;
		rom[ 2337 ] =    -96;
		rom[ 2338 ] =    -67;
		rom[ 2339 ] =     -7;
		rom[ 2340 ] =     52;
		rom[ 2341 ] =    171;
		rom[ 2342 ] =     44;
		rom[ 2343 ] =   -214;
		rom[ 2344 ] =     -8;
		rom[ 2345 ] =    107;
		rom[ 2346 ] =     17;
		rom[ 2347 ] =    -40;
		rom[ 2348 ] =   -181;
		rom[ 2349 ] =    -41;
		rom[ 2350 ] =     99;
		rom[ 2351 ] =      4;
		rom[ 2352 ] =     12;
		rom[ 2353 ] =    -69;
		rom[ 2354 ] =    216;
		rom[ 2355 ] =     39;
		rom[ 2356 ] =   -237;
		rom[ 2357 ] =    132;
		rom[ 2358 ] =     35;
		rom[ 2359 ] =   -230;
		rom[ 2360 ] =     50;
		rom[ 2361 ] =     24;
		rom[ 2362 ] =    -15;
		rom[ 2363 ] =     62;
		rom[ 2364 ] =    156;
		rom[ 2365 ] =    232;
		rom[ 2366 ] =    -80;
		rom[ 2367 ] =   -170;
		rom[ 2368 ] =     15;
		rom[ 2369 ] =    204;
		rom[ 2370 ] =     48;
		rom[ 2371 ] =    150;
		rom[ 2372 ] =    -65;
		rom[ 2373 ] =     -3;
		rom[ 2374 ] =     52;
		rom[ 2375 ] =   -274;
		rom[ 2376 ] =   -148;
		rom[ 2377 ] =   -169;
		rom[ 2378 ] =   -123;
		rom[ 2379 ] =    147;
		rom[ 2380 ] =    -13;
		rom[ 2381 ] =     31;
		rom[ 2382 ] =     28;
		rom[ 2383 ] =   -444;
		rom[ 2384 ] =     34;
		rom[ 2385 ] =   -120;
		rom[ 2386 ] =    178;
		rom[ 2387 ] =    431;
		rom[ 2388 ] =    203;
		rom[ 2389 ] =   -259;
		rom[ 2390 ] =     36;
		rom[ 2391 ] =    129;
		rom[ 2392 ] =    -40;
		rom[ 2393 ] =   -139;
		rom[ 2394 ] =    -44;
		rom[ 2395 ] =     64;
		rom[ 2396 ] =    238;
		rom[ 2397 ] =     -8;
		rom[ 2398 ] =     89;
		rom[ 2399 ] =     17;
		rom[ 2400 ] =     36;
		rom[ 2401 ] =   -263;
		rom[ 2402 ] =    -50;
		rom[ 2403 ] =   -198;
		rom[ 2404 ] =     33;
		rom[ 2405 ] =    -39;
		rom[ 2406 ] =     38;
		rom[ 2407 ] =   -182;
		rom[ 2408 ] =    284;
		rom[ 2409 ] =    238;
		rom[ 2410 ] =    -50;
		rom[ 2411 ] =    107;
		rom[ 2412 ] =   -132;
		rom[ 2413 ] =    -11;
		rom[ 2414 ] =     13;
		rom[ 2415 ] =    -60;
		rom[ 2416 ] =   -226;
		rom[ 2417 ] =    -52;
		rom[ 2418 ] =     34;
		rom[ 2419 ] =    -44;
		rom[ 2420 ] =     14;
		rom[ 2421 ] =     40;
		rom[ 2422 ] =    182;
		rom[ 2423 ] =    -40;
		rom[ 2424 ] =    -88;
		rom[ 2425 ] =   -142;
		rom[ 2426 ] =   -924;
		rom[ 2427 ] =    132;
		rom[ 2428 ] =    -22;
		rom[ 2429 ] =      7;
		rom[ 2430 ] =     60;
		rom[ 2431 ] =    -10;
		rom[ 2432 ] =    117;
		rom[ 2433 ] =   -195;
		rom[ 2434 ] =   -957;
		rom[ 2435 ] =   -163;
		rom[ 2436 ] =     49;
		rom[ 2437 ] =    -41;
		rom[ 2438 ] =      5;
		rom[ 2439 ] =   -434;
		rom[ 2440 ] =    303;
		rom[ 2441 ] =   -104;
		rom[ 2442 ] =     39;
		rom[ 2443 ] =    125;
		rom[ 2444 ] =    -62;
		rom[ 2445 ] =    -12;
		rom[ 2446 ] =    111;
		rom[ 2447 ] =     48;
		rom[ 2448 ] =   -112;
		rom[ 2449 ] =    -52;
		rom[ 2450 ] =     79;
		rom[ 2451 ] =    -79;
		rom[ 2452 ] =     35;
		rom[ 2453 ] =   -130;
		rom[ 2454 ] =    122;
		rom[ 2455 ] =    115;
		rom[ 2456 ] =     33;
		rom[ 2457 ] =    -10;
		rom[ 2458 ] =    -88;
		rom[ 2459 ] =      1;
		rom[ 2460 ] =     20;
		rom[ 2461 ] =    297;
		rom[ 2462 ] =    -82;
		rom[ 2463 ] =    -46;
		rom[ 2464 ] =      0;
		rom[ 2465 ] =    -37;
		rom[ 2466 ] =   -101;
		rom[ 2467 ] =    -46;
		rom[ 2468 ] =     37;
		rom[ 2469 ] =    -15;
		rom[ 2470 ] =     87;
		rom[ 2471 ] =     79;
		rom[ 2472 ] =     -9;
		rom[ 2473 ] =    -45;
		rom[ 2474 ] =   -258;
		rom[ 2475 ] =   -137;
		rom[ 2476 ] =    123;
		rom[ 2477 ] =     67;
		rom[ 2478 ] =      9;
		rom[ 2479 ] =   -153;
		rom[ 2480 ] =     39;
		rom[ 2481 ] =    -37;
		rom[ 2482 ] =      3;
		rom[ 2483 ] =     -4;
		rom[ 2484 ] =     91;
		rom[ 2485 ] =    306;
		rom[ 2486 ] =   -158;
		rom[ 2487 ] =   -467;
		rom[ 2488 ] =  -7680;
		rom[ 2489 ] =    -61;
		rom[ 2490 ] =     -8;
		rom[ 2491 ] =    -39;
		rom[ 2492 ] =    -15;
		rom[ 2493 ] =   -165;
		rom[ 2494 ] =    278;
		rom[ 2495 ] =    -66;
		rom[ 2496 ] =     35;
		rom[ 2497 ] =    -53;
		rom[ 2498 ] =     37;
		rom[ 2499 ] =      7;
		rom[ 2500 ] =    323;
		rom[ 2501 ] =    -32;
		rom[ 2502 ] =   -175;
		rom[ 2503 ] =   -122;
		rom[ 2504 ] =   -120;
		rom[ 2505 ] =     65;
		rom[ 2506 ] =   -123;
		rom[ 2507 ] =    -61;
		rom[ 2508 ] =    194;
		rom[ 2509 ] =    -89;
		rom[ 2510 ] =   -202;
		rom[ 2511 ] =    120;
		rom[ 2512 ] =    171;
		rom[ 2513 ] =     63;
		rom[ 2514 ] =    -55;
		rom[ 2515 ] =     71;
		rom[ 2516 ] =     14;
		rom[ 2517 ] =   -255;
		rom[ 2518 ] =   -305;
		rom[ 2519 ] =     38;
		rom[ 2520 ] =   -363;
		rom[ 2521 ] =    -72;
		rom[ 2522 ] =    121;
		rom[ 2523 ] =    -15;
		rom[ 2524 ] =   -219;
		rom[ 2525 ] =     42;
		rom[ 2526 ] =   -300;
		rom[ 2527 ] =     67;
		rom[ 2528 ] =      9;
		rom[ 2529 ] =    -10;
		rom[ 2530 ] =     73;
		rom[ 2531 ] =   -360;
		rom[ 2532 ] =    -54;
		rom[ 2533 ] =     86;
		rom[ 2534 ] =    -64;
		rom[ 2535 ] =     10;
		rom[ 2536 ] =    135;
		rom[ 2537 ] =     64;
		rom[ 2538 ] =      1;
		rom[ 2539 ] =   -127;
		rom[ 2540 ] =     21;
		rom[ 2541 ] =   -133;
		rom[ 2542 ] =   -161;
		rom[ 2543 ] =    329;
		rom[ 2544 ] =    213;
		rom[ 2545 ] =     28;
		rom[ 2546 ] =   -345;
		rom[ 2547 ] =   -346;
		rom[ 2548 ] =    103;
		rom[ 2549 ] =    -67;
		rom[ 2550 ] =    150;
		rom[ 2551 ] =    -42;
		rom[ 2552 ] =      3;
		rom[ 2553 ] =     -4;
		rom[ 2554 ] =    -61;
		rom[ 2555 ] =   -137;
		rom[ 2556 ] =    192;
		rom[ 2557 ] =    -41;
		rom[ 2558 ] =    -44;
		rom[ 2559 ] =     59;
		rom[ 2560 ] =     64;
		rom[ 2561 ] =     33;
		rom[ 2562 ] =   -214;
		rom[ 2563 ] =    603;
		rom[ 2564 ] =     48;
		rom[ 2565 ] =     37;
		rom[ 2566 ] =    -11;
		rom[ 2567 ] =     45;
		rom[ 2568 ] =   -252;
		rom[ 2569 ] =    -41;
		rom[ 2570 ] =    -61;
		rom[ 2571 ] =     36;
		rom[ 2572 ] =   -266;
		rom[ 2573 ] =     50;
		rom[ 2574 ] =   -232;
		rom[ 2575 ] =     -7;
		rom[ 2576 ] =   -255;
		rom[ 2577 ] =    187;
		rom[ 2578 ] =     71;
		rom[ 2579 ] =      1;
		rom[ 2580 ] =    -51;
		rom[ 2581 ] =    165;
		rom[ 2582 ] =    -47;
		rom[ 2583 ] =    -74;
		rom[ 2584 ] =    -17;
		rom[ 2585 ] =     -3;
		rom[ 2586 ] =    -53;
		rom[ 2587 ] =    -91;
		rom[ 2588 ] =    277;
		rom[ 2589 ] =     54;
		rom[ 2590 ] =    132;
		rom[ 2591 ] =   -112;
		rom[ 2592 ] =      8;
		rom[ 2593 ] =      3;
		rom[ 2594 ] =     87;
		rom[ 2595 ] =     84;
		rom[ 2596 ] =    -64;
		rom[ 2597 ] =     35;
		rom[ 2598 ] =     -3;
		rom[ 2599 ] =     48;
		rom[ 2600 ] =     89;
		rom[ 2601 ] =     -9;
		rom[ 2602 ] =   -109;
		rom[ 2603 ] =    170;
		rom[ 2604 ] =   -125;
		rom[ 2605 ] =     33;
		rom[ 2606 ] =    -14;
		rom[ 2607 ] =   -147;
		rom[ 2608 ] =    249;
		rom[ 2609 ] =     45;
		rom[ 2610 ] =   -207;
		rom[ 2611 ] =     71;
		rom[ 2612 ] =    -34;
		rom[ 2613 ] =    -17;
		rom[ 2614 ] =    -46;
		rom[ 2615 ] =    -40;
		rom[ 2616 ] =     74;
		rom[ 2617 ] =    113;
		rom[ 2618 ] =    -49;
		rom[ 2619 ] =     -2;
		rom[ 2620 ] =   -108;
		rom[ 2621 ] =   -218;
		rom[ 2622 ] =    214;
		rom[ 2623 ] =     25;
		rom[ 2624 ] =    -47;
		rom[ 2625 ] =     64;
		rom[ 2626 ] =    -90;
		rom[ 2627 ] =     41;
		rom[ 2628 ] =    -37;
		rom[ 2629 ] =    -54;
		rom[ 2630 ] =   -182;
		rom[ 2631 ] =      8;
		rom[ 2632 ] =    -69;
		rom[ 2633 ] =     92;
		rom[ 2634 ] =    -12;
		rom[ 2635 ] =     33;
		rom[ 2636 ] =   -275;
		rom[ 2637 ] =      6;
		rom[ 2638 ] =    -66;
		rom[ 2639 ] =   -454;
		rom[ 2640 ] =     76;
		rom[ 2641 ] =     50;
		rom[ 2642 ] =   -110;
		rom[ 2643 ] =   -130;
		rom[ 2644 ] =    199;
		rom[ 2645 ] =   -161;
		rom[ 2646 ] =    -11;
		rom[ 2647 ] =     30;
		rom[ 2648 ] =     -4;
		rom[ 2649 ] =     22;
		rom[ 2650 ] =     10;
		rom[ 2651 ] =   -486;
		rom[ 2652 ] =    -15;
		rom[ 2653 ] =    227;
		rom[ 2654 ] =    -56;
		rom[ 2655 ] =    147;
		rom[ 2656 ] =   -138;
		rom[ 2657 ] =    -20;
		rom[ 2658 ] =    -51;
		rom[ 2659 ] =    106;
		rom[ 2660 ] =     -7;
		rom[ 2661 ] =    -30;
		rom[ 2662 ] =     84;
		rom[ 2663 ] =     -5;
		rom[ 2664 ] =   -112;
		rom[ 2665 ] =     30;
		rom[ 2666 ] =    234;
		rom[ 2667 ] =     28;
		rom[ 2668 ] =    -36;
		rom[ 2669 ] =     51;
		rom[ 2670 ] =     83;
		rom[ 2671 ] =     40;
		rom[ 2672 ] =    -19;
		rom[ 2673 ] =     29;
		rom[ 2674 ] =    -42;
		rom[ 2675 ] =     57;
		rom[ 2676 ] =    -49;
		rom[ 2677 ] =     29;
		rom[ 2678 ] =   -229;
		rom[ 2679 ] =     91;
		rom[ 2680 ] =   -117;
		rom[ 2681 ] =     60;
		rom[ 2682 ] =     -7;
		rom[ 2683 ] =   -130;
		rom[ 2684 ] =   -138;
		rom[ 2685 ] =   -227;
		rom[ 2686 ] =    206;
		rom[ 2687 ] =      3;
		rom[ 2688 ] =    -11;
		rom[ 2689 ] =     18;
		rom[ 2690 ] =    -50;
		rom[ 2691 ] =  -1391;
		rom[ 2692 ] =    114;
		rom[ 2693 ] =     -3;
		rom[ 2694 ] =    -38;
		rom[ 2695 ] =    118;
		rom[ 2696 ] =   -422;
		rom[ 2697 ] =     -9;
		rom[ 2698 ] =     88;
		rom[ 2699 ] =     31;
		rom[ 2700 ] =    -15;
		rom[ 2701 ] =      4;
		rom[ 2702 ] =    -70;
		rom[ 2703 ] =    -45;
		rom[ 2704 ] =    -82;
		rom[ 2705 ] =     32;
		rom[ 2706 ] =   -127;
		rom[ 2707 ] =     11;
		rom[ 2708 ] =    -10;
		rom[ 2709 ] =      0;
		rom[ 2710 ] =   -391;
		rom[ 2711 ] =      9;
		rom[ 2712 ] =     25;
		rom[ 2713 ] =    159;
		rom[ 2714 ] =   -238;
		rom[ 2715 ] =   -103;
		rom[ 2716 ] =     24;
		rom[ 2717 ] =     95;
		rom[ 2718 ] =    -59;
		rom[ 2719 ] =     10;
		rom[ 2720 ] =   -127;
		rom[ 2721 ] =      8;
		rom[ 2722 ] =   -128;
		rom[ 2723 ] =      9;
		rom[ 2724 ] =    -16;
		rom[ 2725 ] =    124;
		rom[ 2726 ] =     34;
		rom[ 2727 ] =   -113;
		rom[ 2728 ] =      7;
		rom[ 2729 ] =      3;
		rom[ 2730 ] =      3;
		rom[ 2731 ] =     74;
		rom[ 2732 ] =   -103;
		rom[ 2733 ] =     84;
		rom[ 2734 ] =   -136;
		rom[ 2735 ] =   -369;
		rom[ 2736 ] =   -202;
		rom[ 2737 ] =    -68;
		rom[ 2738 ] =   -139;
		rom[ 2739 ] =      5;
		rom[ 2740 ] =   -127;
		rom[ 2741 ] =   -202;
		rom[ 2742 ] =    204;
		rom[ 2743 ] =    -84;
		rom[ 2744 ] =    -69;
		rom[ 2745 ] =   -135;
		rom[ 2746 ] =   -144;
		rom[ 2747 ] =    -44;
		rom[ 2748 ] =    -23;
		rom[ 2749 ] =    -14;
		rom[ 2750 ] =     60;
		rom[ 2751 ] =     45;
		rom[ 2752 ] =   -109;
		rom[ 2753 ] =    148;
		rom[ 2754 ] =      8;
		rom[ 2755 ] =     17;
		rom[ 2756 ] =   -321;
		rom[ 2757 ] =    136;
		rom[ 2758 ] =    298;
		rom[ 2759 ] =    100;
		rom[ 2760 ] =   -188;
		rom[ 2761 ] =    -36;
		rom[ 2762 ] =     30;
		rom[ 2763 ] =   -362;
		rom[ 2764 ] =    113;
		rom[ 2765 ] =   -356;
		rom[ 2766 ] =    131;
		rom[ 2767 ] =    -14;
		rom[ 2768 ] =    -20;
		rom[ 2769 ] =   -221;
		rom[ 2770 ] =    133;
		rom[ 2771 ] =    -41;
		rom[ 2772 ] =    -43;
		rom[ 2773 ] =     -1;
		rom[ 2774 ] =    162;
		rom[ 2775 ] =    -86;
		rom[ 2776 ] =     -8;
		rom[ 2777 ] =    165;
		rom[ 2778 ] =     13;
		rom[ 2779 ] =    167;
		rom[ 2780 ] =     49;
		rom[ 2781 ] =   -238;
		rom[ 2782 ] =   -174;
		rom[ 2783 ] =      3;
		rom[ 2784 ] =    257;
		rom[ 2785 ] =    -59;
		rom[ 2786 ] =   -185;
		rom[ 2787 ] =    -56;
		rom[ 2788 ] =     42;
		rom[ 2789 ] =    -61;
		rom[ 2790 ] =    130;
		rom[ 2791 ] =    231;
		rom[ 2792 ] =     35;
		rom[ 2793 ] =   -169;
		rom[ 2794 ] =    205;
		rom[ 2795 ] =    -85;
		rom[ 2796 ] =   -142;
		rom[ 2797 ] =    -15;
		rom[ 2798 ] =     87;
		rom[ 2799 ] =     71;
		rom[ 2800 ] =    300;
		rom[ 2801 ] =    209;
		rom[ 2802 ] =    -47;
		rom[ 2803 ] =     83;
		rom[ 2804 ] =     50;
		rom[ 2805 ] =   -239;
		rom[ 2806 ] =      6;
		rom[ 2807 ] =    -54;
		rom[ 2808 ] =    189;
		rom[ 2809 ] =    -49;
		rom[ 2810 ] =    178;
		rom[ 2811 ] =    100;
		rom[ 2812 ] =    -18;
		rom[ 2813 ] =    244;
		rom[ 2814 ] =    -13;
		rom[ 2815 ] =     19;
		rom[ 2816 ] =     13;
		rom[ 2817 ] =    184;
		rom[ 2818 ] =     36;
		rom[ 2819 ] =     10;
		rom[ 2820 ] =    137;
		rom[ 2821 ] =    -11;
		rom[ 2822 ] =      8;
		rom[ 2823 ] =    -66;
		rom[ 2824 ] =     40;
		rom[ 2825 ] =   -187;
		rom[ 2826 ] =     21;
		rom[ 2827 ] =    -90;
		rom[ 2828 ] =     72;
		rom[ 2829 ] =   -215;
		rom[ 2830 ] =     38;
		rom[ 2831 ] =    -48;
		rom[ 2832 ] =    113;
		rom[ 2833 ] =    -14;
		rom[ 2834 ] =    -79;
		rom[ 2835 ] =    420;
		rom[ 2836 ] =   -199;
		rom[ 2837 ] =    -59;
		rom[ 2838 ] =    -92;
		rom[ 2839 ] =    199;
		rom[ 2840 ] =    302;
		rom[ 2841 ] =   -120;
		rom[ 2842 ] =     56;
		rom[ 2843 ] =     -9;
		rom[ 2844 ] =    107;
		rom[ 2845 ] =    -42;
		rom[ 2846 ] =     40;
		rom[ 2847 ] =     -1;
		rom[ 2848 ] =     -7;
		rom[ 2849 ] =    -58;
		rom[ 2850 ] =    -15;
		rom[ 2851 ] =    -76;
		rom[ 2852 ] =     56;
		rom[ 2853 ] =    311;
		rom[ 2854 ] =      3;
		rom[ 2855 ] =   -382;
		rom[ 2856 ] =    -98;
		rom[ 2857 ] =    -54;
		rom[ 2858 ] =      0;
		rom[ 2859 ] =   -159;
		rom[ 2860 ] =   -108;
		rom[ 2861 ] =      6;
		rom[ 2862 ] =     33;
		rom[ 2863 ] =    301;
		rom[ 2864 ] =      8;
		rom[ 2865 ] =    -81;
		rom[ 2866 ] =    216;
		rom[ 2867 ] =     94;
		rom[ 2868 ] =   -133;
		rom[ 2869 ] =    -15;
		rom[ 2870 ] =    202;
		rom[ 2871 ] =   -299;
		rom[ 2872 ] =     10;
		rom[ 2873 ] =    -91;
		rom[ 2874 ] =     53;
		rom[ 2875 ] =    -48;
		rom[ 2876 ] =     65;
		rom[ 2877 ] =      8;
		rom[ 2878 ] =   -253;
		rom[ 2879 ] =    -34;
		rom[ 2880 ] =     86;
		rom[ 2881 ] =    -46;
		rom[ 2882 ] =   -251;
		rom[ 2883 ] =     -8;
		rom[ 2884 ] =    298;
		rom[ 2885 ] =    163;
		rom[ 2886 ] =    -59;
		rom[ 2887 ] =    -56;
		rom[ 2888 ] =     41;
		rom[ 2889 ] =    -43;
		rom[ 2890 ] =     66;
		rom[ 2891 ] =   -196;
		rom[ 2892 ] =    -69;
		rom[ 2893 ] =     19;
		rom[ 2894 ] =     -9;
		rom[ 2895 ] =    -45;
		rom[ 2896 ] =     48;
		rom[ 2897 ] =    180;
		rom[ 2898 ] =     17;
		rom[ 2899 ] =    192;
		rom[ 2900 ] =     49;
		rom[ 2901 ] =    -12;
		rom[ 2902 ] =   -114;
		rom[ 2903 ] =    166;
		rom[ 2904 ] =    -14;
		rom[ 2905 ] =    -39;
		rom[ 2906 ] =   -156;
		rom[ 2907 ] =    -12;
		rom[ 2908 ] =     28;
		rom[ 2909 ] =   -204;
		rom[ 2910 ] =    -48;
		rom[ 2911 ] =    -34;
		rom[ 2912 ] =    124;
	end
endmodule

module right_tree_rom(
	input 				clk,
	input		[11:0]	addr,
	output reg	[13:0]	q    // x y w h 5bit*4
	);
	reg					[13:0]	rom [4095:0];
	always @(posedge clk) q <= rom[addr];
	initial begin
		rom[ 0    ] =   -567;
		rom[ 1    ] =    339;
		rom[ 2    ] =    272;
		rom[ 3    ] =    301;
		rom[ 4    ] =    322;
		rom[ 5    ] =   -479;
		rom[ 6    ] =    112;
		rom[ 7    ] =    113;
		rom[ 8    ] =    218;
		rom[ 9    ] =   -402;
		rom[ 10   ] =    302;
		rom[ 11   ] =    179;
		rom[ 12   ] =    442;
		rom[ 13   ] =   -558;
		rom[ 14   ] =    116;
		rom[ 15   ] =    137;
		rom[ 16   ] =    238;
		rom[ 17   ] =   -169;
		rom[ 18   ] =    -76;
		rom[ 19   ] =    347;
		rom[ 20   ] =    -50;
		rom[ 21   ] =   -135;
		rom[ 22   ] =    292;
		rom[ 23   ] =    197;
		rom[ 24   ] =   -387;
		rom[ 25   ] =    375;
		rom[ 26   ] =    256;
		rom[ 27   ] =   -408;
		rom[ 28   ] =    212;
		rom[ 29   ] =    108;
		rom[ 30   ] =    269;
		rom[ 31   ] =   -344;
		rom[ 32   ] =    371;
		rom[ 33   ] =    310;
		rom[ 34   ] =   -117;
		rom[ 35   ] =     39;
		rom[ 36   ] =   -400;
		rom[ 37   ] =     59;
		rom[ 38   ] =    327;
		rom[ 39   ] =    -77;
		rom[ 40   ] =    -13;
		rom[ 41   ] =    393;
		rom[ 42   ] =    239;
		rom[ 43   ] =    246;
		rom[ 44   ] =   -757;
		rom[ 45   ] =   -112;
		rom[ 46   ] =    102;
		rom[ 47   ] =   -677;
		rom[ 48   ] =     72;
		rom[ 49   ] =     59;
		rom[ 50   ] =    275;
		rom[ 51   ] =     25;
		rom[ 52   ] =   -274;
		rom[ 53   ] =    196;
		rom[ 54   ] =    353;
		rom[ 55   ] =    132;
		rom[ 56   ] =    149;
		rom[ 57   ] =    299;
		rom[ 58   ] =    244;
		rom[ 59   ] =    -35;
		rom[ 60   ] =     70;
		rom[ 61   ] =     60;
		rom[ 62   ] =   -343;
		rom[ 63   ] =   -230;
		rom[ 64   ] =   -418;
		rom[ 65   ] =     46;
		rom[ 66   ] =    -97;
		rom[ 67   ] =     63;
		rom[ 68   ] =    -75;
		rom[ 69   ] =    161;
		rom[ 70   ] =     13;
		rom[ 71   ] =     99;
		rom[ 72   ] =     25;
		rom[ 73   ] =   -322;
		rom[ 74   ] =   -609;
		rom[ 75   ] =    -70;
		rom[ 76   ] =   -291;
		rom[ 77   ] =   -324;
		rom[ 78   ] =     69;
		rom[ 79   ] =    181;
		rom[ 80   ] =      9;
		rom[ 81   ] =    -12;
		rom[ 82   ] =    -89;
		rom[ 83   ] =     54;
		rom[ 84   ] =    277;
		rom[ 85   ] =    359;
		rom[ 86   ] =    189;
		rom[ 87   ] =     96;
		rom[ 88   ] =    323;
		rom[ 89   ] =    117;
		rom[ 90   ] =   -245;
		rom[ 91   ] =     11;
		rom[ 92   ] =    138;
		rom[ 93   ] =   -381;
		rom[ 94   ] =   -134;
		rom[ 95   ] =   -409;
		rom[ 96   ] =     39;
		rom[ 97   ] =   -184;
		rom[ 98   ] =     17;
		rom[ 99   ] =    174;
		rom[ 100  ] =     19;
		rom[ 101  ] =    -55;
		rom[ 102  ] =    335;
		rom[ 103  ] =    312;
		rom[ 104  ] =    217;
		rom[ 105  ] =     76;
		rom[ 106  ] =    -83;
		rom[ 107  ] =   -214;
		rom[ 108  ] =   -171;
		rom[ 109  ] =     35;
		rom[ 110  ] =     19;
		rom[ 111  ] =     49;
		rom[ 112  ] =     17;
		rom[ 113  ] =    199;
		rom[ 114  ] =     31;
		rom[ 115  ] =      3;
		rom[ 116  ] =    135;
		rom[ 117  ] =    100;
		rom[ 118  ] =   -542;
		rom[ 119  ] =    252;
		rom[ 120  ] =     24;
		rom[ 121  ] =    -37;
		rom[ 122  ] =   -148;
		rom[ 123  ] =    -43;
		rom[ 124  ] =   -163;
		rom[ 125  ] =     64;
		rom[ 126  ] =    -69;
		rom[ 127  ] =     60;
		rom[ 128  ] =   -323;
		rom[ 129  ] =     77;
		rom[ 130  ] =    135;
		rom[ 131  ] =     61;
		rom[ 132  ] =    132;
		rom[ 133  ] =     -3;
		rom[ 134  ] =    -66;
		rom[ 135  ] =   -151;
		rom[ 136  ] =    267;
		rom[ 137  ] =    141;
		rom[ 138  ] =    163;
		rom[ 139  ] =    136;
		rom[ 140  ] =     92;
		rom[ 141  ] =     92;
		rom[ 142  ] =   -128;
		rom[ 143  ] =    218;
		rom[ 144  ] =    292;
		rom[ 145  ] =    -46;
		rom[ 146  ] =    -80;
		rom[ 147  ] =    267;
		rom[ 148  ] =     50;
		rom[ 149  ] =   -340;
		rom[ 150  ] =   -179;
		rom[ 151  ] =     57;
		rom[ 152  ] =   -131;
		rom[ 153  ] =    158;
		rom[ 154  ] =    121;
		rom[ 155  ] =   -175;
		rom[ 156  ] =     29;
		rom[ 157  ] =    -14;
		rom[ 158  ] =    211;
		rom[ 159  ] =    -45;
		rom[ 160  ] =   -396;
		rom[ 161  ] =     61;
		rom[ 162  ] =    -81;
		rom[ 163  ] =   -211;
		rom[ 164  ] =     13;
		rom[ 165  ] =     33;
		rom[ 166  ] =      9;
		rom[ 167  ] =    126;
		rom[ 168  ] =   -146;
		rom[ 169  ] =    163;
		rom[ 170  ] =     16;
		rom[ 171  ] =   -255;
		rom[ 172  ] =      9;
		rom[ 173  ] =   -266;
		rom[ 174  ] =   -138;
		rom[ 175  ] =    113;
		rom[ 176  ] =      0;
		rom[ 177  ] =   -165;
		rom[ 178  ] =    205;
		rom[ 179  ] =     54;
		rom[ 180  ] =   -270;
		rom[ 181  ] =   -219;
		rom[ 182  ] =     16;
		rom[ 183  ] =    162;
		rom[ 184  ] =    144;
		rom[ 185  ] =   -385;
		rom[ 186  ] =     96;
		rom[ 187  ] =     31;
		rom[ 188  ] =    173;
		rom[ 189  ] =    243;
		rom[ 190  ] =    125;
		rom[ 191  ] =    127;
		rom[ 192  ] =   -320;
		rom[ 193  ] =    152;
		rom[ 194  ] =     77;
		rom[ 195  ] =     57;
		rom[ 196  ] =    -25;
		rom[ 197  ] =     47;
		rom[ 198  ] =   -119;
		rom[ 199  ] =    -67;
		rom[ 200  ] =    106;
		rom[ 201  ] =    151;
		rom[ 202  ] =   -117;
		rom[ 203  ] =     36;
		rom[ 204  ] =   -249;
		rom[ 205  ] =     46;
		rom[ 206  ] =   -339;
		rom[ 207  ] =   -536;
		rom[ 208  ] =    131;
		rom[ 209  ] =   -328;
		rom[ 210  ] =   -118;
		rom[ 211  ] =     11;
		rom[ 212  ] =     88;
		rom[ 213  ] =    109;
		rom[ 214  ] =     42;
		rom[ 215  ] =   -120;
		rom[ 216  ] =   -427;
		rom[ 217  ] =      9;
		rom[ 218  ] =     59;
		rom[ 219  ] =     25;
		rom[ 220  ] =    -48;
		rom[ 221  ] =    -97;
		rom[ 222  ] =     50;
		rom[ 223  ] =    129;
		rom[ 224  ] =     59;
		rom[ 225  ] =    -81;
		rom[ 226  ] =     -3;
		rom[ 227  ] =    266;
		rom[ 228  ] =   -213;
		rom[ 229  ] =    116;
		rom[ 230  ] =   -384;
		rom[ 231  ] =    -98;
		rom[ 232  ] =    -27;
		rom[ 233  ] =   -430;
		rom[ 234  ] =     61;
		rom[ 235  ] =    119;
		rom[ 236  ] =     45;
		rom[ 237  ] =     18;
		rom[ 238  ] =   -395;
		rom[ 239  ] =     96;
		rom[ 240  ] =   -317;
		rom[ 241  ] =     13;
		rom[ 242  ] =     58;
		rom[ 243  ] =    314;
		rom[ 244  ] =    -11;
		rom[ 245  ] =    -55;
		rom[ 246  ] =   -486;
		rom[ 247  ] =      1;
		rom[ 248  ] =    -21;
		rom[ 249  ] =     16;
		rom[ 250  ] =   -195;
		rom[ 251  ] =    210;
		rom[ 252  ] =     75;
		rom[ 253  ] =    148;
		rom[ 254  ] =    229;
		rom[ 255  ] =    129;
		rom[ 256  ] =   -180;
		rom[ 257  ] =    181;
		rom[ 258  ] =     68;
		rom[ 259  ] =    -98;
		rom[ 260  ] =     66;
		rom[ 261  ] =   -150;
		rom[ 262  ] =     43;
		rom[ 263  ] =   -224;
		rom[ 264  ] =     60;
		rom[ 265  ] =   -144;
		rom[ 266  ] =     98;
		rom[ 267  ] =   -355;
		rom[ 268  ] =   -273;
		rom[ 269  ] =     50;
		rom[ 270  ] =    111;
		rom[ 271  ] =   -114;
		rom[ 272  ] =     57;
		rom[ 273  ] =     -1;
		rom[ 274  ] =   -133;
		rom[ 275  ] =   -386;
		rom[ 276  ] =     47;
		rom[ 277  ] =      0;
		rom[ 278  ] =   -568;
		rom[ 279  ] =     15;
		rom[ 280  ] =   -303;
		rom[ 281  ] =     31;
		rom[ 282  ] =    181;
		rom[ 283  ] =   -269;
		rom[ 284  ] =     49;
		rom[ 285  ] =    -64;
		rom[ 286  ] =    -54;
		rom[ 287  ] =    -71;
		rom[ 288  ] =     62;
		rom[ 289  ] =     14;
		rom[ 290  ] =     50;
		rom[ 291  ] =    269;
		rom[ 292  ] =   -440;
		rom[ 293  ] =     15;
		rom[ 294  ] =      7;
		rom[ 295  ] =   -123;
		rom[ 296  ] =     41;
		rom[ 297  ] =     10;
		rom[ 298  ] =     82;
		rom[ 299  ] =    -67;
		rom[ 300  ] =     38;
		rom[ 301  ] =     10;
		rom[ 302  ] =     39;
		rom[ 303  ] =   -108;
		rom[ 304  ] =     47;
		rom[ 305  ] =      0;
		rom[ 306  ] =     79;
		rom[ 307  ] =   -166;
		rom[ 308  ] =     39;
		rom[ 309  ] =    391;
		rom[ 310  ] =    166;
		rom[ 311  ] =      9;
		rom[ 312  ] =    -25;
		rom[ 313  ] =    -87;
		rom[ 314  ] =     -4;
		rom[ 315  ] =     -7;
		rom[ 316  ] =     42;
		rom[ 317  ] =      0;
		rom[ 318  ] =    -45;
		rom[ 319  ] =   -327;
		rom[ 320  ] =   -388;
		rom[ 321  ] =     83;
		rom[ 322  ] =     38;
		rom[ 323  ] =    284;
		rom[ 324  ] =   -157;
		rom[ 325  ] =    101;
		rom[ 326  ] =     73;
		rom[ 327  ] =    115;
		rom[ 328  ] =   -174;
		rom[ 329  ] =     15;
		rom[ 330  ] =   -442;
		rom[ 331  ] =     31;
		rom[ 332  ] =   -207;
		rom[ 333  ] =    172;
		rom[ 334  ] =    215;
		rom[ 335  ] =   -121;
		rom[ 336  ] =    242;
		rom[ 337  ] =    -80;
		rom[ 338  ] =     45;
		rom[ 339  ] =     63;
		rom[ 340  ] =   -109;
		rom[ 341  ] =   -409;
		rom[ 342  ] =     96;
		rom[ 343  ] =     63;
		rom[ 344  ] =   -369;
		rom[ 345  ] =   -348;
		rom[ 346  ] =     69;
		rom[ 347  ] =   -208;
		rom[ 348  ] =   -191;
		rom[ 349  ] =    207;
		rom[ 350  ] =    220;
		rom[ 351  ] =   -253;
		rom[ 352  ] =     39;
		rom[ 353  ] =   -180;
		rom[ 354  ] =   -103;
		rom[ 355  ] =     18;
		rom[ 356  ] =   -184;
		rom[ 357  ] =     67;
		rom[ 358  ] =     37;
		rom[ 359  ] =   -275;
		rom[ 360  ] =    311;
		rom[ 361  ] =      3;
		rom[ 362  ] =    -39;
		rom[ 363  ] =    180;
		rom[ 364  ] =     85;
		rom[ 365  ] =     19;
		rom[ 366  ] =     12;
		rom[ 367  ] =    -62;
		rom[ 368  ] =     31;
		rom[ 369  ] =     -6;
		rom[ 370  ] =    -30;
		rom[ 371  ] =    -68;
		rom[ 372  ] =   -165;
		rom[ 373  ] =   -317;
		rom[ 374  ] =    260;
		rom[ 375  ] =    -92;
		rom[ 376  ] =     52;
		rom[ 377  ] =     -5;
		rom[ 378  ] =    -75;
		rom[ 379  ] =    277;
		rom[ 380  ] =    311;
		rom[ 381  ] =   -272;
		rom[ 382  ] =     43;
		rom[ 383  ] =    132;
		rom[ 384  ] =     63;
		rom[ 385  ] =   -592;
		rom[ 386  ] =    -83;
		rom[ 387  ] =     18;
		rom[ 388  ] =   -441;
		rom[ 389  ] =    260;
		rom[ 390  ] =     38;
		rom[ 391  ] =    -74;
		rom[ 392  ] =    -86;
		rom[ 393  ] =   -600;
		rom[ 394  ] =     39;
		rom[ 395  ] =     -7;
		rom[ 396  ] =     60;
		rom[ 397  ] =    236;
		rom[ 398  ] =     79;
		rom[ 399  ] =   -693;
		rom[ 400  ] =     -8;
		rom[ 401  ] =     58;
		rom[ 402  ] =   -267;
		rom[ 403  ] =    196;
		rom[ 404  ] =     71;
		rom[ 405  ] =    -65;
		rom[ 406  ] =    280;
		rom[ 407  ] =    135;
		rom[ 408  ] =    103;
		rom[ 409  ] =    189;
		rom[ 410  ] =    188;
		rom[ 411  ] =     97;
		rom[ 412  ] =     93;
		rom[ 413  ] =    203;
		rom[ 414  ] =    -84;
		rom[ 415  ] =   -247;
		rom[ 416  ] =   -271;
		rom[ 417  ] =     34;
		rom[ 418  ] =    154;
		rom[ 419  ] =    -54;
		rom[ 420  ] =   -375;
		rom[ 421  ] =     52;
		rom[ 422  ] =     26;
		rom[ 423  ] =   -102;
		rom[ 424  ] =   -411;
		rom[ 425  ] =    -34;
		rom[ 426  ] =      2;
		rom[ 427  ] =     66;
		rom[ 428  ] =   -183;
		rom[ 429  ] =   -421;
		rom[ 430  ] =      6;
		rom[ 431  ] =    -26;
		rom[ 432  ] =   -137;
		rom[ 433  ] =     51;
		rom[ 434  ] =   -258;
		rom[ 435  ] =    -70;
		rom[ 436  ] =   -136;
		rom[ 437  ] =     53;
		rom[ 438  ] =     -9;
		rom[ 439  ] =   -182;
		rom[ 440  ] =      4;
		rom[ 441  ] =    -16;
		rom[ 442  ] =    203;
		rom[ 443  ] =   -175;
		rom[ 444  ] =    -55;
		rom[ 445  ] =    319;
		rom[ 446  ] =     37;
		rom[ 447  ] =     -3;
		rom[ 448  ] =    276;
		rom[ 449  ] =    291;
		rom[ 450  ] =     -1;
		rom[ 451  ] =     61;
		rom[ 452  ] =    -52;
		rom[ 453  ] =   -312;
		rom[ 454  ] =     13;
		rom[ 455  ] =     74;
		rom[ 456  ] =   -171;
		rom[ 457  ] =      4;
		rom[ 458  ] =      6;
		rom[ 459  ] =      7;
		rom[ 460  ] =    151;
		rom[ 461  ] =     67;
		rom[ 462  ] =    -85;
		rom[ 463  ] =     40;
		rom[ 464  ] =     -6;
		rom[ 465  ] =    -11;
		rom[ 466  ] =   -114;
		rom[ 467  ] =     36;
		rom[ 468  ] =    -97;
		rom[ 469  ] =     16;
		rom[ 470  ] =    203;
		rom[ 471  ] =     29;
		rom[ 472  ] =     -1;
		rom[ 473  ] =    104;
		rom[ 474  ] =    -98;
		rom[ 475  ] =    196;
		rom[ 476  ] =    -57;
		rom[ 477  ] =   -372;
		rom[ 478  ] =     66;
		rom[ 479  ] =    124;
		rom[ 480  ] =    -56;
		rom[ 481  ] =     37;
		rom[ 482  ] =    -51;
		rom[ 483  ] =     69;
		rom[ 484  ] =    -48;
		rom[ 485  ] =     40;
		rom[ 486  ] =   -419;
		rom[ 487  ] =     61;
		rom[ 488  ] =     -1;
		rom[ 489  ] =   -115;
		rom[ 490  ] =    112;
		rom[ 491  ] =     64;
		rom[ 492  ] =      6;
		rom[ 493  ] =      0;
		rom[ 494  ] =    389;
		rom[ 495  ] =    -55;
		rom[ 496  ] =      5;
		rom[ 497  ] =    164;
		rom[ 498  ] =    147;
		rom[ 499  ] =    336;
		rom[ 500  ] =     74;
		rom[ 501  ] =    136;
		rom[ 502  ] =   -114;
		rom[ 503  ] =    -70;
		rom[ 504  ] =     52;
		rom[ 505  ] =     17;
		rom[ 506  ] =   -133;
		rom[ 507  ] =     11;
		rom[ 508  ] =     47;
		rom[ 509  ] =   -176;
		rom[ 510  ] =   -215;
		rom[ 511  ] =   -349;
		rom[ 512  ] =     66;
		rom[ 513  ] =     16;
		rom[ 514  ] =     -4;
		rom[ 515  ] =    -83;
		rom[ 516  ] =     51;
		rom[ 517  ] =     57;
		rom[ 518  ] =   -274;
		rom[ 519  ] =      9;
		rom[ 520  ] =   -183;
		rom[ 521  ] =   -136;
		rom[ 522  ] =    249;
		rom[ 523  ] =    -60;
		rom[ 524  ] =    117;
		rom[ 525  ] =   -682;
		rom[ 526  ] =      6;
		rom[ 527  ] =   -555;
		rom[ 528  ] =    191;
		rom[ 529  ] =      2;
		rom[ 530  ] =    254;
		rom[ 531  ] =    -63;
		rom[ 532  ] =   -156;
		rom[ 533  ] =      7;
		rom[ 534  ] =    -34;
		rom[ 535  ] =   -133;
		rom[ 536  ] =     38;
		rom[ 537  ] =      0;
		rom[ 538  ] =   -157;
		rom[ 539  ] =    -53;
		rom[ 540  ] =    122;
		rom[ 541  ] =     28;
		rom[ 542  ] =   -383;
		rom[ 543  ] =    208;
		rom[ 544  ] =    -17;
		rom[ 545  ] =     12;
		rom[ 546  ] =     -1;
		rom[ 547  ] =    -47;
		rom[ 548  ] =     24;
		rom[ 549  ] =    -69;
		rom[ 550  ] =     40;
		rom[ 551  ] =    -60;
		rom[ 552  ] =     50;
		rom[ 553  ] =      5;
		rom[ 554  ] =     -4;
		rom[ 555  ] =   -444;
		rom[ 556  ] =    -14;
		rom[ 557  ] =   -197;
		rom[ 558  ] =    171;
		rom[ 559  ] =     79;
		rom[ 560  ] =     65;
		rom[ 561  ] =    105;
		rom[ 562  ] =      4;
		rom[ 563  ] =    -53;
		rom[ 564  ] =     10;
		rom[ 565  ] =     43;
		rom[ 566  ] =    209;
		rom[ 567  ] =      6;
		rom[ 568  ] =    -87;
		rom[ 569  ] =      0;
		rom[ 570  ] =     64;
		rom[ 571  ] =   -366;
		rom[ 572  ] =     85;
		rom[ 573  ] =     33;
		rom[ 574  ] =    -79;
		rom[ 575  ] =    181;
		rom[ 576  ] =     49;
		rom[ 577  ] =   -227;
		rom[ 578  ] =    -70;
		rom[ 579  ] =      6;
		rom[ 580  ] =    -44;
		rom[ 581  ] =    -51;
		rom[ 582  ] =     29;
		rom[ 583  ] =   -116;
		rom[ 584  ] =    100;
		rom[ 585  ] =    -51;
		rom[ 586  ] =     52;
		rom[ 587  ] =   -261;
		rom[ 588  ] =    -23;
		rom[ 589  ] =   -493;
		rom[ 590  ] =    -17;
		rom[ 591  ] =     47;
		rom[ 592  ] =     56;
		rom[ 593  ] =    -47;
		rom[ 594  ] =     95;
		rom[ 595  ] =    -68;
		rom[ 596  ] =    147;
		rom[ 597  ] =    258;
		rom[ 598  ] =    144;
		rom[ 599  ] =     79;
		rom[ 600  ] =   -286;
		rom[ 601  ] =     84;
		rom[ 602  ] =    134;
		rom[ 603  ] =     -8;
		rom[ 604  ] =     30;
		rom[ 605  ] =     53;
		rom[ 606  ] =    -72;
		rom[ 607  ] =   -179;
		rom[ 608  ] =    187;
		rom[ 609  ] =     39;
		rom[ 610  ] =    -87;
		rom[ 611  ] =    -33;
		rom[ 612  ] =   -245;
		rom[ 613  ] =   -119;
		rom[ 614  ] =   -134;
		rom[ 615  ] =     55;
		rom[ 616  ] =     16;
		rom[ 617  ] =     55;
		rom[ 618  ] =     12;
		rom[ 619  ] =     44;
		rom[ 620  ] =    -56;
		rom[ 621  ] =     46;
		rom[ 622  ] =     14;
		rom[ 623  ] =    134;
		rom[ 624  ] =    143;
		rom[ 625  ] =   -179;
		rom[ 626  ] =     11;
		rom[ 627  ] =     66;
		rom[ 628  ] =    148;
		rom[ 629  ] =     50;
		rom[ 630  ] =     54;
		rom[ 631  ] =    197;
		rom[ 632  ] =    -63;
		rom[ 633  ] =     -9;
		rom[ 634  ] =    282;
		rom[ 635  ] =    184;
		rom[ 636  ] =     11;
		rom[ 637  ] =    -96;
		rom[ 638  ] =    286;
		rom[ 639  ] =     49;
		rom[ 640  ] =   -297;
		rom[ 641  ] =     42;
		rom[ 642  ] =     -3;
		rom[ 643  ] =    -21;
		rom[ 644  ] =    152;
		rom[ 645  ] =     34;
		rom[ 646  ] =     -8;
		rom[ 647  ] =      4;
		rom[ 648  ] =    136;
		rom[ 649  ] =     41;
		rom[ 650  ] =   -192;
		rom[ 651  ] =   -167;
		rom[ 652  ] =   -314;
		rom[ 653  ] =    110;
		rom[ 654  ] =   -305;
		rom[ 655  ] =     36;
		rom[ 656  ] =    138;
		rom[ 657  ] =    144;
		rom[ 658  ] =   -203;
		rom[ 659  ] =    379;
		rom[ 660  ] =     -7;
		rom[ 661  ] =      8;
		rom[ 662  ] =     76;
		rom[ 663  ] =    -97;
		rom[ 664  ] =   -135;
		rom[ 665  ] =    538;
		rom[ 666  ] =    -10;
		rom[ 667  ] =     91;
		rom[ 668  ] =    -45;
		rom[ 669  ] =   -332;
		rom[ 670  ] =     35;
		rom[ 671  ] =    100;
		rom[ 672  ] =   -184;
		rom[ 673  ] =     16;
		rom[ 674  ] =    -42;
		rom[ 675  ] =    -42;
		rom[ 676  ] =    187;
		rom[ 677  ] =     52;
		rom[ 678  ] =    -75;
		rom[ 679  ] =    103;
		rom[ 680  ] =    -44;
		rom[ 681  ] =    178;
		rom[ 682  ] =      0;
		rom[ 683  ] =    137;
		rom[ 684  ] =   -191;
		rom[ 685  ] =     85;
		rom[ 686  ] =     -9;
		rom[ 687  ] =      4;
		rom[ 688  ] =    186;
		rom[ 689  ] =   -125;
		rom[ 690  ] =    197;
		rom[ 691  ] =     17;
		rom[ 692  ] =    -47;
		rom[ 693  ] =   -410;
		rom[ 694  ] =    304;
		rom[ 695  ] =    100;
		rom[ 696  ] =   -412;
		rom[ 697  ] =    138;
		rom[ 698  ] =    -81;
		rom[ 699  ] =   -263;
		rom[ 700  ] =   -202;
		rom[ 701  ] =   -214;
		rom[ 702  ] =   -160;
		rom[ 703  ] =    402;
		rom[ 704  ] =     98;
		rom[ 705  ] =    134;
		rom[ 706  ] =    -72;
		rom[ 707  ] =    -78;
		rom[ 708  ] =   -223;
		rom[ 709  ] =    -51;
		rom[ 710  ] =     20;
		rom[ 711  ] =    145;
		rom[ 712  ] =    114;
		rom[ 713  ] =    173;
		rom[ 714  ] =     49;
		rom[ 715  ] =   -182;
		rom[ 716  ] =     29;
		rom[ 717  ] =     51;
		rom[ 718  ] =     93;
		rom[ 719  ] =     32;
		rom[ 720  ] =    147;
		rom[ 721  ] =   -134;
		rom[ 722  ] =    122;
		rom[ 723  ] =   -398;
		rom[ 724  ] =     48;
		rom[ 725  ] =   -114;
		rom[ 726  ] =    -54;
		rom[ 727  ] =    133;
		rom[ 728  ] =      7;
		rom[ 729  ] =    -57;
		rom[ 730  ] =     37;
		rom[ 731  ] =      4;
		rom[ 732  ] =   -252;
		rom[ 733  ] =      5;
		rom[ 734  ] =     50;
		rom[ 735  ] =     97;
		rom[ 736  ] =    -37;
		rom[ 737  ] =    -71;
		rom[ 738  ] =    154;
		rom[ 739  ] =    -96;
		rom[ 740  ] =    264;
		rom[ 741  ] =    -57;
		rom[ 742  ] =   -303;
		rom[ 743  ] =     11;
		rom[ 744  ] =    274;
		rom[ 745  ] =    -44;
		rom[ 746  ] =    -18;
		rom[ 747  ] =    102;
		rom[ 748  ] =   -311;
		rom[ 749  ] =   -182;
		rom[ 750  ] =     46;
		rom[ 751  ] =   -395;
		rom[ 752  ] =     42;
		rom[ 753  ] =     -4;
		rom[ 754  ] =     60;
		rom[ 755  ] =     14;
		rom[ 756  ] =     -4;
		rom[ 757  ] =    -54;
		rom[ 758  ] =     47;
		rom[ 759  ] =   -101;
		rom[ 760  ] =   -657;
		rom[ 761  ] =     -3;
		rom[ 762  ] =     42;
		rom[ 763  ] =     84;
		rom[ 764  ] =   -124;
		rom[ 765  ] =    -57;
		rom[ 766  ] =     48;
		rom[ 767  ] =    -53;
		rom[ 768  ] =   -153;
		rom[ 769  ] =     -5;
		rom[ 770  ] =     15;
		rom[ 771  ] =   -394;
		rom[ 772  ] =     95;
		rom[ 773  ] =     35;
		rom[ 774  ] =     -4;
		rom[ 775  ] =   -313;
		rom[ 776  ] =      0;
		rom[ 777  ] =     -3;
		rom[ 778  ] =   -317;
		rom[ 779  ] =    131;
		rom[ 780  ] =   -181;
		rom[ 781  ] =      0;
		rom[ 782  ] =     37;
		rom[ 783  ] =   -119;
		rom[ 784  ] =   -106;
		rom[ 785  ] =    111;
		rom[ 786  ] =   -243;
		rom[ 787  ] =    -78;
		rom[ 788  ] =   -506;
		rom[ 789  ] =     -2;
		rom[ 790  ] =     -8;
		rom[ 791  ] =     99;
		rom[ 792  ] =    150;
		rom[ 793  ] =   -242;
		rom[ 794  ] =     54;
		rom[ 795  ] =     -7;
		rom[ 796  ] =    297;
		rom[ 797  ] =   -285;
		rom[ 798  ] =     53;
		rom[ 799  ] =    -40;
		rom[ 800  ] =     46;
		rom[ 801  ] =     11;
		rom[ 802  ] =   -191;
		rom[ 803  ] =   -428;
		rom[ 804  ] =    195;
		rom[ 805  ] =   -226;
		rom[ 806  ] =   -630;
		rom[ 807  ] =    -76;
		rom[ 808  ] =     41;
		rom[ 809  ] =    -95;
		rom[ 810  ] =    152;
		rom[ 811  ] =    141;
		rom[ 812  ] =    104;
		rom[ 813  ] =    -60;
		rom[ 814  ] =     40;
		rom[ 815  ] =    -87;
		rom[ 816  ] =     24;
		rom[ 817  ] =      8;
		rom[ 818  ] =    -13;
		rom[ 819  ] =     -5;
		rom[ 820  ] =    234;
		rom[ 821  ] =    -73;
		rom[ 822  ] =    136;
		rom[ 823  ] =   -113;
		rom[ 824  ] =   -655;
		rom[ 825  ] =   -283;
		rom[ 826  ] =    145;
		rom[ 827  ] =     32;
		rom[ 828  ] =    223;
		rom[ 829  ] =     53;
		rom[ 830  ] =     14;
		rom[ 831  ] =     -2;
		rom[ 832  ] =     43;
		rom[ 833  ] =   -355;
		rom[ 834  ] =      0;
		rom[ 835  ] =   -106;
		rom[ 836  ] =      4;
		rom[ 837  ] =    -50;
		rom[ 838  ] =    132;
		rom[ 839  ] =    180;
		rom[ 840  ] =   -171;
		rom[ 841  ] =     91;
		rom[ 842  ] =     48;
		rom[ 843  ] =     67;
		rom[ 844  ] =     68;
		rom[ 845  ] =   -276;
		rom[ 846  ] =    -71;
		rom[ 847  ] =     61;
		rom[ 848  ] =    -63;
		rom[ 849  ] =      1;
		rom[ 850  ] =    181;
		rom[ 851  ] =   -368;
		rom[ 852  ] =     12;
		rom[ 853  ] =   -114;
		rom[ 854  ] =     88;
		rom[ 855  ] =   -343;
		rom[ 856  ] =   -132;
		rom[ 857  ] =   -186;
		rom[ 858  ] =     -6;
		rom[ 859  ] =     49;
		rom[ 860  ] =   -224;
		rom[ 861  ] =    -61;
		rom[ 862  ] =   -320;
		rom[ 863  ] =    -21;
		rom[ 864  ] =   -124;
		rom[ 865  ] =     46;
		rom[ 866  ] =    159;
		rom[ 867  ] =    236;
		rom[ 868  ] =    198;
		rom[ 869  ] =   -278;
		rom[ 870  ] =    -59;
		rom[ 871  ] =    158;
		rom[ 872  ] =    258;
		rom[ 873  ] =     11;
		rom[ 874  ] =      1;
		rom[ 875  ] =      4;
		rom[ 876  ] =    -73;
		rom[ 877  ] =    -42;
		rom[ 878  ] =     -2;
		rom[ 879  ] =    -75;
		rom[ 880  ] =     -7;
		rom[ 881  ] =   -182;
		rom[ 882  ] =   -388;
		rom[ 883  ] =    -99;
		rom[ 884  ] =     -5;
		rom[ 885  ] =     37;
		rom[ 886  ] =   -105;
		rom[ 887  ] =    105;
		rom[ 888  ] =    141;
		rom[ 889  ] =      4;
		rom[ 890  ] =    -75;
		rom[ 891  ] =   -118;
		rom[ 892  ] =   -132;
		rom[ 893  ] =     53;
		rom[ 894  ] =    367;
		rom[ 895  ] =    -10;
		rom[ 896  ] =     34;
		rom[ 897  ] =     27;
		rom[ 898  ] =     57;
		rom[ 899  ] =     96;
		rom[ 900  ] =    -50;
		rom[ 901  ] =    149;
		rom[ 902  ] =   -171;
		rom[ 903  ] =    -19;
		rom[ 904  ] =    298;
		rom[ 905  ] =     11;
		rom[ 906  ] =    -55;
		rom[ 907  ] =     51;
		rom[ 908  ] =     10;
		rom[ 909  ] =     91;
		rom[ 910  ] =     49;
		rom[ 911  ] =     62;
		rom[ 912  ] =    325;
		rom[ 913  ] =   -551;
		rom[ 914  ] =    -41;
		rom[ 915  ] =     54;
		rom[ 916  ] =    -50;
		rom[ 917  ] =     55;
		rom[ 918  ] =   -255;
		rom[ 919  ] =    125;
		rom[ 920  ] =    -44;
		rom[ 921  ] =   -191;
		rom[ 922  ] =    139;
		rom[ 923  ] =   -129;
		rom[ 924  ] =   -245;
		rom[ 925  ] =     43;
		rom[ 926  ] =   -336;
		rom[ 927  ] =      3;
		rom[ 928  ] =     61;
		rom[ 929  ] =     39;
		rom[ 930  ] =     -3;
		rom[ 931  ] =     16;
		rom[ 932  ] =    -11;
		rom[ 933  ] =     39;
		rom[ 934  ] =     13;
		rom[ 935  ] =      1;
		rom[ 936  ] =   -341;
		rom[ 937  ] =     95;
		rom[ 938  ] =    -38;
		rom[ 939  ] =     65;
		rom[ 940  ] =   -267;
		rom[ 941  ] =    101;
		rom[ 942  ] =      8;
		rom[ 943  ] =     96;
		rom[ 944  ] =    -53;
		rom[ 945  ] =     45;
		rom[ 946  ] =   -165;
		rom[ 947  ] =   -253;
		rom[ 948  ] =      8;
		rom[ 949  ] =      0;
		rom[ 950  ] =    120;
		rom[ 951  ] =    146;
		rom[ 952  ] =   -487;
		rom[ 953  ] =     -2;
		rom[ 954  ] =    -13;
		rom[ 955  ] =   -314;
		rom[ 956  ] =   -277;
		rom[ 957  ] =    -94;
		rom[ 958  ] =     60;
		rom[ 959  ] =     39;
		rom[ 960  ] =   -486;
		rom[ 961  ] =      5;
		rom[ 962  ] =    156;
		rom[ 963  ] =     47;
		rom[ 964  ] =    550;
		rom[ 965  ] =     33;
		rom[ 966  ] =   -132;
		rom[ 967  ] =    316;
		rom[ 968  ] =     -8;
		rom[ 969  ] =    411;
		rom[ 970  ] =     -1;
		rom[ 971  ] =    243;
		rom[ 972  ] =    495;
		rom[ 973  ] =   -178;
		rom[ 974  ] =     78;
		rom[ 975  ] =    146;
		rom[ 976  ] =    148;
		rom[ 977  ] =    110;
		rom[ 978  ] =    -51;
		rom[ 979  ] =    281;
		rom[ 980  ] =     14;
		rom[ 981  ] =    -85;
		rom[ 982  ] =     57;
		rom[ 983  ] =     15;
		rom[ 984  ] =     47;
		rom[ 985  ] =    -66;
		rom[ 986  ] =    182;
		rom[ 987  ] =     19;
		rom[ 988  ] =    232;
		rom[ 989  ] =    185;
		rom[ 990  ] =     53;
		rom[ 991  ] =     -3;
		rom[ 992  ] =    -29;
		rom[ 993  ] =   -196;
		rom[ 994  ] =     10;
		rom[ 995  ] =    151;
		rom[ 996  ] =     83;
		rom[ 997  ] =    -65;
		rom[ 998  ] =   -143;
		rom[ 999  ] =   -134;
		rom[ 1000 ] =     75;
		rom[ 1001 ] =     64;
		rom[ 1002 ] =   -120;
		rom[ 1003 ] =   -289;
		rom[ 1004 ] =    -67;
		rom[ 1005 ] =     -4;
		rom[ 1006 ] =     40;
		rom[ 1007 ] =   -179;
		rom[ 1008 ] =     59;
		rom[ 1009 ] =    116;
		rom[ 1010 ] =     36;
		rom[ 1011 ] =    -65;
		rom[ 1012 ] =   -453;
		rom[ 1013 ] =    138;
		rom[ 1014 ] =     85;
		rom[ 1015 ] =   -298;
		rom[ 1016 ] =   -638;
		rom[ 1017 ] =    245;
		rom[ 1018 ] =    -65;
		rom[ 1019 ] =   -258;
		rom[ 1020 ] =     49;
		rom[ 1021 ] =   -256;
		rom[ 1022 ] =    106;
		rom[ 1023 ] =    100;
		rom[ 1024 ] =    -92;
		rom[ 1025 ] =    237;
		rom[ 1026 ] =     85;
		rom[ 1027 ] =     23;
		rom[ 1028 ] =     62;
		rom[ 1029 ] =   -322;
		rom[ 1030 ] =     43;
		rom[ 1031 ] =   -224;
		rom[ 1032 ] =     33;
		rom[ 1033 ] =     56;
		rom[ 1034 ] =   -129;
		rom[ 1035 ] =    117;
		rom[ 1036 ] =    142;
		rom[ 1037 ] =      4;
		rom[ 1038 ] =    -43;
		rom[ 1039 ] =      1;
		rom[ 1040 ] =     28;
		rom[ 1041 ] =    -47;
		rom[ 1042 ] =    210;
		rom[ 1043 ] =    -88;
		rom[ 1044 ] =   -356;
		rom[ 1045 ] =      0;
		rom[ 1046 ] =     29;
		rom[ 1047 ] =     -6;
		rom[ 1048 ] =     30;
		rom[ 1049 ] =    -53;
		rom[ 1050 ] =    136;
		rom[ 1051 ] =    -79;
		rom[ 1052 ] =    -13;
		rom[ 1053 ] =     -3;
		rom[ 1054 ] =    107;
		rom[ 1055 ] =     10;
		rom[ 1056 ] =    162;
		rom[ 1057 ] =      2;
		rom[ 1058 ] =    -16;
		rom[ 1059 ] =     21;
		rom[ 1060 ] =   -102;
		rom[ 1061 ] =    131;
		rom[ 1062 ] =     35;
		rom[ 1063 ] =    160;
		rom[ 1064 ] =   -698;
		rom[ 1065 ] =   -276;
		rom[ 1066 ] =      8;
		rom[ 1067 ] =    112;
		rom[ 1068 ] =    -61;
		rom[ 1069 ] =    -78;
		rom[ 1070 ] =     66;
		rom[ 1071 ] =   -501;
		rom[ 1072 ] =    189;
		rom[ 1073 ] =     67;
		rom[ 1074 ] =     43;
		rom[ 1075 ] =    -66;
		rom[ 1076 ] =    -73;
		rom[ 1077 ] =   -451;
		rom[ 1078 ] =     -6;
		rom[ 1079 ] =    263;
		rom[ 1080 ] =   -319;
		rom[ 1081 ] =   -439;
		rom[ 1082 ] =     52;
		rom[ 1083 ] =     52;
		rom[ 1084 ] =     51;
		rom[ 1085 ] =    427;
		rom[ 1086 ] =    -90;
		rom[ 1087 ] =    -46;
		rom[ 1088 ] =     31;
		rom[ 1089 ] =   -296;
		rom[ 1090 ] =  -1198;
		rom[ 1091 ] =    -37;
		rom[ 1092 ] =     87;
		rom[ 1093 ] =     78;
		rom[ 1094 ] =      6;
		rom[ 1095 ] =     55;
		rom[ 1096 ] =     40;
		rom[ 1097 ] =     -2;
		rom[ 1098 ] =   -176;
		rom[ 1099 ] =    311;
		rom[ 1100 ] =   -105;
		rom[ 1101 ] =     -4;
		rom[ 1102 ] =     49;
		rom[ 1103 ] =   -107;
		rom[ 1104 ] =    200;
		rom[ 1105 ] =     -8;
		rom[ 1106 ] =     16;
		rom[ 1107 ] =    -48;
		rom[ 1108 ] =   -202;
		rom[ 1109 ] =    150;
		rom[ 1110 ] =    -75;
		rom[ 1111 ] =    106;
		rom[ 1112 ] =     43;
		rom[ 1113 ] =      6;
		rom[ 1114 ] =   -106;
		rom[ 1115 ] =     91;
		rom[ 1116 ] =    220;
		rom[ 1117 ] =     25;
		rom[ 1118 ] =   -177;
		rom[ 1119 ] =      9;
		rom[ 1120 ] =   -177;
		rom[ 1121 ] =   -247;
		rom[ 1122 ] =      0;
		rom[ 1123 ] =    -83;
		rom[ 1124 ] =    185;
		rom[ 1125 ] =     77;
		rom[ 1126 ] =    -26;
		rom[ 1127 ] =    -55;
		rom[ 1128 ] =    -40;
		rom[ 1129 ] =     -5;
		rom[ 1130 ] =    -97;
		rom[ 1131 ] =    -69;
		rom[ 1132 ] =     67;
		rom[ 1133 ] =    142;
		rom[ 1134 ] =      7;
		rom[ 1135 ] =     16;
		rom[ 1136 ] =    -53;
		rom[ 1137 ] =     16;
		rom[ 1138 ] =     71;
		rom[ 1139 ] =   -226;
		rom[ 1140 ] =     40;
		rom[ 1141 ] =    108;
		rom[ 1142 ] =     40;
		rom[ 1143 ] =     31;
		rom[ 1144 ] =    210;
		rom[ 1145 ] =    -43;
		rom[ 1146 ] =     37;
		rom[ 1147 ] =     -7;
		rom[ 1148 ] =   -177;
		rom[ 1149 ] =     -6;
		rom[ 1150 ] =     37;
		rom[ 1151 ] =      9;
		rom[ 1152 ] =    205;
		rom[ 1153 ] =    -63;
		rom[ 1154 ] =     50;
		rom[ 1155 ] =     34;
		rom[ 1156 ] =     47;
		rom[ 1157 ] =    -89;
		rom[ 1158 ] =     53;
		rom[ 1159 ] =     -3;
		rom[ 1160 ] =   -116;
		rom[ 1161 ] =      3;
		rom[ 1162 ] =      8;
		rom[ 1163 ] =     69;
		rom[ 1164 ] =     44;
		rom[ 1165 ] =     17;
		rom[ 1166 ] =     30;
		rom[ 1167 ] =    284;
		rom[ 1168 ] =    117;
		rom[ 1169 ] =    -47;
		rom[ 1170 ] =     36;
		rom[ 1171 ] =      2;
		rom[ 1172 ] =   -282;
		rom[ 1173 ] =      0;
		rom[ 1174 ] =     89;
		rom[ 1175 ] =     -7;
		rom[ 1176 ] =    -37;
		rom[ 1177 ] =   -634;
		rom[ 1178 ] =   -112;
		rom[ 1179 ] =    180;
		rom[ 1180 ] =    157;
		rom[ 1181 ] =     -6;
		rom[ 1182 ] =   -275;
		rom[ 1183 ] =   -181;
		rom[ 1184 ] =      8;
		rom[ 1185 ] =     44;
		rom[ 1186 ] =      3;
		rom[ 1187 ] =    287;
		rom[ 1188 ] =     44;
		rom[ 1189 ] =    -46;
		rom[ 1190 ] =    -61;
		rom[ 1191 ] =      0;
		rom[ 1192 ] =     66;
		rom[ 1193 ] =     66;
		rom[ 1194 ] =    150;
		rom[ 1195 ] =    -55;
		rom[ 1196 ] =     39;
		rom[ 1197 ] =   -290;
		rom[ 1198 ] =    318;
		rom[ 1199 ] =    -48;
		rom[ 1200 ] =     31;
		rom[ 1201 ] =      2;
		rom[ 1202 ] =    -29;
		rom[ 1203 ] =    -14;
		rom[ 1204 ] =    -10;
		rom[ 1205 ] =   -276;
		rom[ 1206 ] =      0;
		rom[ 1207 ] =   -216;
		rom[ 1208 ] =   -203;
		rom[ 1209 ] =    -54;
		rom[ 1210 ] =    109;
		rom[ 1211 ] =      0;
		rom[ 1212 ] =     57;
		rom[ 1213 ] =    -98;
		rom[ 1214 ] =   -203;
		rom[ 1215 ] =    104;
		rom[ 1216 ] =    203;
		rom[ 1217 ] =     29;
		rom[ 1218 ] =    320;
		rom[ 1219 ] =    197;
		rom[ 1220 ] =     40;
		rom[ 1221 ] =   -471;
		rom[ 1222 ] =    -39;
		rom[ 1223 ] =      0;
		rom[ 1224 ] =     43;
		rom[ 1225 ] =      1;
		rom[ 1226 ] =     63;
		rom[ 1227 ] =   -469;
		rom[ 1228 ] =    -98;
		rom[ 1229 ] =      5;
		rom[ 1230 ] =     -3;
		rom[ 1231 ] =    -72;
		rom[ 1232 ] =   -360;
		rom[ 1233 ] =    204;
		rom[ 1234 ] =    -21;
		rom[ 1235 ] =    -56;
		rom[ 1236 ] =   -330;
		rom[ 1237 ] =    139;
		rom[ 1238 ] =    -41;
		rom[ 1239 ] =    136;
		rom[ 1240 ] =    -43;
		rom[ 1241 ] =     10;
		rom[ 1242 ] =   -264;
		rom[ 1243 ] =     81;
		rom[ 1244 ] =   -418;
		rom[ 1245 ] =    -51;
		rom[ 1246 ] =   -172;
		rom[ 1247 ] =    231;
		rom[ 1248 ] =   -327;
		rom[ 1249 ] =    193;
		rom[ 1250 ] =     57;
		rom[ 1251 ] =     79;
		rom[ 1252 ] =    -98;
		rom[ 1253 ] =     70;
		rom[ 1254 ] =   -310;
		rom[ 1255 ] =    -79;
		rom[ 1256 ] =    -52;
		rom[ 1257 ] =     52;
		rom[ 1258 ] =      9;
		rom[ 1259 ] =     40;
		rom[ 1260 ] =    302;
		rom[ 1261 ] =     84;
		rom[ 1262 ] =    106;
		rom[ 1263 ] =     45;
		rom[ 1264 ] =   -114;
		rom[ 1265 ] =    -28;
		rom[ 1266 ] =    -10;
		rom[ 1267 ] =    -12;
		rom[ 1268 ] =    -52;
		rom[ 1269 ] =   -290;
		rom[ 1270 ] =      4;
		rom[ 1271 ] =     57;
		rom[ 1272 ] =     10;
		rom[ 1273 ] =   -285;
		rom[ 1274 ] =    -37;
		rom[ 1275 ] =  -1014;
		rom[ 1276 ] =   -252;
		rom[ 1277 ] =   -191;
		rom[ 1278 ] =     77;
		rom[ 1279 ] =    134;
		rom[ 1280 ] =     -1;
		rom[ 1281 ] =     60;
		rom[ 1282 ] =     20;
		rom[ 1283 ] =   -171;
		rom[ 1284 ] =    -53;
		rom[ 1285 ] =   -267;
		rom[ 1286 ] =      0;
		rom[ 1287 ] =    157;
		rom[ 1288 ] =   -217;
		rom[ 1289 ] =   -130;
		rom[ 1290 ] =   -325;
		rom[ 1291 ] =    696;
		rom[ 1292 ] =     39;
		rom[ 1293 ] =     35;
		rom[ 1294 ] =     87;
		rom[ 1295 ] =    123;
		rom[ 1296 ] =   -514;
		rom[ 1297 ] =    -28;
		rom[ 1298 ] =   -298;
		rom[ 1299 ] =     36;
		rom[ 1300 ] =    157;
		rom[ 1301 ] =   -192;
		rom[ 1302 ] =    256;
		rom[ 1303 ] =     -8;
		rom[ 1304 ] =    -47;
		rom[ 1305 ] =     74;
		rom[ 1306 ] =    152;
		rom[ 1307 ] =     45;
		rom[ 1308 ] =    -54;
		rom[ 1309 ] =    154;
		rom[ 1310 ] =     -6;
		rom[ 1311 ] =    145;
		rom[ 1312 ] =    -69;
		rom[ 1313 ] =     63;
		rom[ 1314 ] =    -52;
		rom[ 1315 ] =   -194;
		rom[ 1316 ] =    -65;
		rom[ 1317 ] =    -73;
		rom[ 1318 ] =      8;
		rom[ 1319 ] =    -68;
		rom[ 1320 ] =   -293;
		rom[ 1321 ] =     76;
		rom[ 1322 ] =   -339;
		rom[ 1323 ] =    180;
		rom[ 1324 ] =   -115;
		rom[ 1325 ] =    -15;
		rom[ 1326 ] =    112;
		rom[ 1327 ] =    180;
		rom[ 1328 ] =     61;
		rom[ 1329 ] =     29;
		rom[ 1330 ] =   -280;
		rom[ 1331 ] =     19;
		rom[ 1332 ] =     29;
		rom[ 1333 ] =     42;
		rom[ 1334 ] =   -218;
		rom[ 1335 ] =    107;
		rom[ 1336 ] =   -166;
		rom[ 1337 ] =     39;
		rom[ 1338 ] =    -87;
		rom[ 1339 ] =    202;
		rom[ 1340 ] =    -57;
		rom[ 1341 ] =     -1;
		rom[ 1342 ] =    -15;
		rom[ 1343 ] =     51;
		rom[ 1344 ] =    -57;
		rom[ 1345 ] =     63;
		rom[ 1346 ] =    186;
		rom[ 1347 ] =     73;
		rom[ 1348 ] =   -285;
		rom[ 1349 ] =    170;
		rom[ 1350 ] =    -67;
		rom[ 1351 ] =     48;
		rom[ 1352 ] =   -281;
		rom[ 1353 ] =   -750;
		rom[ 1354 ] =    -70;
		rom[ 1355 ] =   -160;
		rom[ 1356 ] =    -94;
		rom[ 1357 ] =     49;
		rom[ 1358 ] =   -498;
		rom[ 1359 ] =     47;
		rom[ 1360 ] =    -39;
		rom[ 1361 ] =     28;
		rom[ 1362 ] =      5;
		rom[ 1363 ] =    252;
		rom[ 1364 ] =    -11;
		rom[ 1365 ] =   -301;
		rom[ 1366 ] =   -239;
		rom[ 1367 ] =   -383;
		rom[ 1368 ] =    400;
		rom[ 1369 ] =   -173;
		rom[ 1370 ] =     27;
		rom[ 1371 ] =      7;
		rom[ 1372 ] =    -43;
		rom[ 1373 ] =     33;
		rom[ 1374 ] =   -133;
		rom[ 1375 ] =     33;
		rom[ 1376 ] =    124;
		rom[ 1377 ] =      2;
		rom[ 1378 ] =    138;
		rom[ 1379 ] =     -5;
		rom[ 1380 ] =    127;
		rom[ 1381 ] =    -56;
		rom[ 1382 ] =      4;
		rom[ 1383 ] =     18;
		rom[ 1384 ] =     -2;
		rom[ 1385 ] =    -73;
		rom[ 1386 ] =   -571;
		rom[ 1387 ] =    104;
		rom[ 1388 ] =    -51;
		rom[ 1389 ] =     69;
		rom[ 1390 ] =     22;
		rom[ 1391 ] =   -280;
		rom[ 1392 ] =    -37;
		rom[ 1393 ] =   -108;
		rom[ 1394 ] =    -52;
		rom[ 1395 ] =      7;
		rom[ 1396 ] =    -55;
		rom[ 1397 ] =     36;
		rom[ 1398 ] =     -3;
		rom[ 1399 ] =     32;
		rom[ 1400 ] =   -162;
		rom[ 1401 ] =   -120;
		rom[ 1402 ] =    499;
		rom[ 1403 ] =   -542;
		rom[ 1404 ] =    126;
		rom[ 1405 ] =    195;
		rom[ 1406 ] =    101;
		rom[ 1407 ] =   -162;
		rom[ 1408 ] =   -147;
		rom[ 1409 ] =   -175;
		rom[ 1410 ] =     70;
		rom[ 1411 ] =     62;
		rom[ 1412 ] =     69;
		rom[ 1413 ] =     29;
		rom[ 1414 ] =     61;
		rom[ 1415 ] =   -169;
		rom[ 1416 ] =    107;
		rom[ 1417 ] =    -48;
		rom[ 1418 ] =   -234;
		rom[ 1419 ] =    100;
		rom[ 1420 ] =    113;
		rom[ 1421 ] =      0;
		rom[ 1422 ] =     43;
		rom[ 1423 ] =   -205;
		rom[ 1424 ] =     46;
		rom[ 1425 ] =    -53;
		rom[ 1426 ] =     56;
		rom[ 1427 ] =    -48;
		rom[ 1428 ] =     37;
		rom[ 1429 ] =    -60;
		rom[ 1430 ] =     55;
		rom[ 1431 ] =   -154;
		rom[ 1432 ] =     39;
		rom[ 1433 ] =      3;
		rom[ 1434 ] =    -23;
		rom[ 1435 ] =   -358;
		rom[ 1436 ] =   -126;
		rom[ 1437 ] =     -3;
		rom[ 1438 ] =      0;
		rom[ 1439 ] =    -75;
		rom[ 1440 ] =     51;
		rom[ 1441 ] =     12;
		rom[ 1442 ] =     38;
		rom[ 1443 ] =    -67;
		rom[ 1444 ] =    266;
		rom[ 1445 ] =   -301;
		rom[ 1446 ] =    -14;
		rom[ 1447 ] =    -62;
		rom[ 1448 ] =     43;
		rom[ 1449 ] =   -273;
		rom[ 1450 ] =   -342;
		rom[ 1451 ] =    116;
		rom[ 1452 ] =    -95;
		rom[ 1453 ] =      4;
		rom[ 1454 ] =     60;
		rom[ 1455 ] =    -82;
		rom[ 1456 ] =   -261;
		rom[ 1457 ] =    -44;
		rom[ 1458 ] =     61;
		rom[ 1459 ] =    -53;
		rom[ 1460 ] =     44;
		rom[ 1461 ] =     -8;
		rom[ 1462 ] =    257;
		rom[ 1463 ] =   -153;
		rom[ 1464 ] =     96;
		rom[ 1465 ] =   -183;
		rom[ 1466 ] =     82;
		rom[ 1467 ] =   -198;
		rom[ 1468 ] =    -15;
		rom[ 1469 ] =    147;
		rom[ 1470 ] =     32;
		rom[ 1471 ] =    -13;
		rom[ 1472 ] =   -162;
		rom[ 1473 ] =    -46;
		rom[ 1474 ] =   -543;
		rom[ 1475 ] =     22;
		rom[ 1476 ] =      4;
		rom[ 1477 ] =   -282;
		rom[ 1478 ] =    -98;
		rom[ 1479 ] =    -43;
		rom[ 1480 ] =    -98;
		rom[ 1481 ] =     90;
		rom[ 1482 ] =   -233;
		rom[ 1483 ] =     -5;
		rom[ 1484 ] =      0;
		rom[ 1485 ] =     88;
		rom[ 1486 ] =     89;
		rom[ 1487 ] =     10;
		rom[ 1488 ] =    -13;
		rom[ 1489 ] =    -82;
		rom[ 1490 ] =   2560;
		rom[ 1491 ] =     85;
		rom[ 1492 ] =     45;
		rom[ 1493 ] =     42;
		rom[ 1494 ] =   -394;
		rom[ 1495 ] =   -255;
		rom[ 1496 ] =      3;
		rom[ 1497 ] =    -51;
		rom[ 1498 ] =    277;
		rom[ 1499 ] =     50;
		rom[ 1500 ] =     17;
		rom[ 1501 ] =   -215;
		rom[ 1502 ] =     93;
		rom[ 1503 ] =    -70;
		rom[ 1504 ] =     27;
		rom[ 1505 ] =    -59;
		rom[ 1506 ] =     44;
		rom[ 1507 ] =   -214;
		rom[ 1508 ] =    -44;
		rom[ 1509 ] =    -37;
		rom[ 1510 ] =      3;
		rom[ 1511 ] =   -194;
		rom[ 1512 ] =    195;
		rom[ 1513 ] =     -2;
		rom[ 1514 ] =     56;
		rom[ 1515 ] =    -91;
		rom[ 1516 ] =     66;
		rom[ 1517 ] =      7;
		rom[ 1518 ] =   -171;
		rom[ 1519 ] =    -37;
		rom[ 1520 ] =     53;
		rom[ 1521 ] =     12;
		rom[ 1522 ] =     33;
		rom[ 1523 ] =    102;
		rom[ 1524 ] =   -182;
		rom[ 1525 ] =    -74;
		rom[ 1526 ] =      0;
		rom[ 1527 ] =     -2;
		rom[ 1528 ] =   -301;
		rom[ 1529 ] =   -475;
		rom[ 1530 ] =     99;
		rom[ 1531 ] =   -284;
		rom[ 1532 ] =    252;
		rom[ 1533 ] =   -177;
		rom[ 1534 ] =     17;
		rom[ 1535 ] =   -639;
		rom[ 1536 ] =     38;
		rom[ 1537 ] =   -547;
		rom[ 1538 ] =    200;
		rom[ 1539 ] =   -184;
		rom[ 1540 ] =   -349;
		rom[ 1541 ] =    186;
		rom[ 1542 ] =     49;
		rom[ 1543 ] =    -10;
		rom[ 1544 ] =      0;
		rom[ 1545 ] =   -465;
		rom[ 1546 ] =     53;
		rom[ 1547 ] =   -362;
		rom[ 1548 ] =    -30;
		rom[ 1549 ] =     66;
		rom[ 1550 ] =     44;
		rom[ 1551 ] =   -156;
		rom[ 1552 ] =     77;
		rom[ 1553 ] =    -58;
		rom[ 1554 ] =     53;
		rom[ 1555 ] =     17;
		rom[ 1556 ] =    133;
		rom[ 1557 ] =   -126;
		rom[ 1558 ] =     20;
		rom[ 1559 ] =    128;
		rom[ 1560 ] =   -149;
		rom[ 1561 ] =    153;
		rom[ 1562 ] =     55;
		rom[ 1563 ] =    156;
		rom[ 1564 ] =    129;
		rom[ 1565 ] =    105;
		rom[ 1566 ] =     24;
		rom[ 1567 ] =     60;
		rom[ 1568 ] =     46;
		rom[ 1569 ] =     10;
		rom[ 1570 ] =   -209;
		rom[ 1571 ] =     57;
		rom[ 1572 ] =    -50;
		rom[ 1573 ] =    206;
		rom[ 1574 ] =      5;
		rom[ 1575 ] =    -19;
		rom[ 1576 ] =    108;
		rom[ 1577 ] =     39;
		rom[ 1578 ] =      2;
		rom[ 1579 ] =   -232;
		rom[ 1580 ] =    -66;
		rom[ 1581 ] =     68;
		rom[ 1582 ] =     25;
		rom[ 1583 ] =     57;
		rom[ 1584 ] =    -67;
		rom[ 1585 ] =     35;
		rom[ 1586 ] =   -185;
		rom[ 1587 ] =    131;
		rom[ 1588 ] =   -277;
		rom[ 1589 ] =     37;
		rom[ 1590 ] =      7;
		rom[ 1591 ] =     64;
		rom[ 1592 ] =    119;
		rom[ 1593 ] =     33;
		rom[ 1594 ] =    -61;
		rom[ 1595 ] =   -157;
		rom[ 1596 ] =      8;
		rom[ 1597 ] =     44;
		rom[ 1598 ] =    -70;
		rom[ 1599 ] =     61;
		rom[ 1600 ] =     36;
		rom[ 1601 ] =    -61;
		rom[ 1602 ] =   -242;
		rom[ 1603 ] =     24;
		rom[ 1604 ] =   -220;
		rom[ 1605 ] =     98;
		rom[ 1606 ] =      7;
		rom[ 1607 ] =     12;
		rom[ 1608 ] =    -61;
		rom[ 1609 ] =     64;
		rom[ 1610 ] =    -59;
		rom[ 1611 ] =    -52;
		rom[ 1612 ] =    -10;
		rom[ 1613 ] =    154;
		rom[ 1614 ] =    229;
		rom[ 1615 ] =    -69;
		rom[ 1616 ] =      5;
		rom[ 1617 ] =    163;
		rom[ 1618 ] =    -59;
		rom[ 1619 ] =      8;
		rom[ 1620 ] =      8;
		rom[ 1621 ] =     42;
		rom[ 1622 ] =   -508;
		rom[ 1623 ] =     97;
		rom[ 1624 ] =   -235;
		rom[ 1625 ] =     58;
		rom[ 1626 ] =    138;
		rom[ 1627 ] =    -32;
		rom[ 1628 ] =     82;
		rom[ 1629 ] =   -155;
		rom[ 1630 ] =     -7;
		rom[ 1631 ] =      7;
		rom[ 1632 ] =    -11;
		rom[ 1633 ] =      2;
		rom[ 1634 ] =    -38;
		rom[ 1635 ] =     43;
		rom[ 1636 ] =    121;
		rom[ 1637 ] =    -89;
		rom[ 1638 ] =    -10;
		rom[ 1639 ] =     40;
		rom[ 1640 ] =    -51;
		rom[ 1641 ] =     22;
		rom[ 1642 ] =     -1;
		rom[ 1643 ] =     36;
		rom[ 1644 ] =      1;
		rom[ 1645 ] =     38;
		rom[ 1646 ] =   -115;
		rom[ 1647 ] =     71;
		rom[ 1648 ] =    172;
		rom[ 1649 ] =     23;
		rom[ 1650 ] =     85;
		rom[ 1651 ] =     35;
		rom[ 1652 ] =   -174;
		rom[ 1653 ] =    138;
		rom[ 1654 ] =    201;
		rom[ 1655 ] =   -122;
		rom[ 1656 ] =   -156;
		rom[ 1657 ] =    106;
		rom[ 1658 ] =    189;
		rom[ 1659 ] =    -34;
		rom[ 1660 ] =    157;
		rom[ 1661 ] =     37;
		rom[ 1662 ] =   -279;
		rom[ 1663 ] =     57;
		rom[ 1664 ] =     14;
		rom[ 1665 ] =    -54;
		rom[ 1666 ] =    158;
		rom[ 1667 ] =     64;
		rom[ 1668 ] =     10;
		rom[ 1669 ] =      0;
		rom[ 1670 ] =    -86;
		rom[ 1671 ] =      2;
		rom[ 1672 ] =    123;
		rom[ 1673 ] =    -44;
		rom[ 1674 ] =      2;
		rom[ 1675 ] =     81;
		rom[ 1676 ] =    -44;
		rom[ 1677 ] =     -2;
		rom[ 1678 ] =    121;
		rom[ 1679 ] =    -68;
		rom[ 1680 ] =   -261;
		rom[ 1681 ] =    146;
		rom[ 1682 ] =   -107;
		rom[ 1683 ] =    737;
		rom[ 1684 ] =    534;
		rom[ 1685 ] =     36;
		rom[ 1686 ] =    138;
		rom[ 1687 ] =   -400;
		rom[ 1688 ] =    -37;
		rom[ 1689 ] =     33;
		rom[ 1690 ] =    -14;
		rom[ 1691 ] =    147;
		rom[ 1692 ] =      5;
		rom[ 1693 ] =     95;
		rom[ 1694 ] =    -58;
		rom[ 1695 ] =   -104;
		rom[ 1696 ] =   -433;
		rom[ 1697 ] =   -117;
		rom[ 1698 ] =     39;
		rom[ 1699 ] =      8;
		rom[ 1700 ] =    -47;
		rom[ 1701 ] =   -122;
		rom[ 1702 ] =    -67;
		rom[ 1703 ] =     13;
		rom[ 1704 ] =    -34;
		rom[ 1705 ] =   -173;
		rom[ 1706 ] =   -187;
		rom[ 1707 ] =     78;
		rom[ 1708 ] =     -8;
		rom[ 1709 ] =     83;
		rom[ 1710 ] =    111;
		rom[ 1711 ] =  -1218;
		rom[ 1712 ] =    -15;
		rom[ 1713 ] =     -8;
		rom[ 1714 ] =   -196;
		rom[ 1715 ] =    -21;
		rom[ 1716 ] =     -6;
		rom[ 1717 ] =   -570;
		rom[ 1718 ] =    -61;
		rom[ 1719 ] =     32;
		rom[ 1720 ] =    -50;
		rom[ 1721 ] =     35;
		rom[ 1722 ] =      7;
		rom[ 1723 ] =    -36;
		rom[ 1724 ] =    -12;
		rom[ 1725 ] =    -17;
		rom[ 1726 ] =    -10;
		rom[ 1727 ] =    209;
		rom[ 1728 ] =    -48;
		rom[ 1729 ] =    155;
		rom[ 1730 ] =    112;
		rom[ 1731 ] =    140;
		rom[ 1732 ] =    118;
		rom[ 1733 ] =   -251;
		rom[ 1734 ] =    182;
		rom[ 1735 ] =    -55;
		rom[ 1736 ] =     64;
		rom[ 1737 ] =   -276;
		rom[ 1738 ] =    131;
		rom[ 1739 ] =   -318;
		rom[ 1740 ] =     52;
		rom[ 1741 ] =    -89;
		rom[ 1742 ] =     52;
		rom[ 1743 ] =      5;
		rom[ 1744 ] =    140;
		rom[ 1745 ] =     68;
		rom[ 1746 ] =   -261;
		rom[ 1747 ] =   -223;
		rom[ 1748 ] =    205;
		rom[ 1749 ] =     58;
		rom[ 1750 ] =     36;
		rom[ 1751 ] =   -489;
		rom[ 1752 ] =    -83;
		rom[ 1753 ] =      0;
		rom[ 1754 ] =     42;
		rom[ 1755 ] =    213;
		rom[ 1756 ] =    -18;
		rom[ 1757 ] =   -295;
		rom[ 1758 ] =     38;
		rom[ 1759 ] =    129;
		rom[ 1760 ] =     74;
		rom[ 1761 ] =   -228;
		rom[ 1762 ] =    -11;
		rom[ 1763 ] =     -5;
		rom[ 1764 ] =    247;
		rom[ 1765 ] =    -44;
		rom[ 1766 ] =     70;
		rom[ 1767 ] =   -455;
		rom[ 1768 ] =     -6;
		rom[ 1769 ] =   -180;
		rom[ 1770 ] =     84;
		rom[ 1771 ] =    -77;
		rom[ 1772 ] =    148;
		rom[ 1773 ] =     11;
		rom[ 1774 ] =     48;
		rom[ 1775 ] =   -176;
		rom[ 1776 ] =     39;
		rom[ 1777 ] =   -153;
		rom[ 1778 ] =     96;
		rom[ 1779 ] =    132;
		rom[ 1780 ] =     36;
		rom[ 1781 ] =    302;
		rom[ 1782 ] =    234;
		rom[ 1783 ] =    -14;
		rom[ 1784 ] =   -256;
		rom[ 1785 ] =     -1;
		rom[ 1786 ] =   -431;
		rom[ 1787 ] =    -39;
		rom[ 1788 ] =    -47;
		rom[ 1789 ] =     -4;
		rom[ 1790 ] =    -65;
		rom[ 1791 ] =    -79;
		rom[ 1792 ] =    107;
		rom[ 1793 ] =    237;
		rom[ 1794 ] =    103;
		rom[ 1795 ] =   -253;
		rom[ 1796 ] =     65;
		rom[ 1797 ] =     30;
		rom[ 1798 ] =   -263;
		rom[ 1799 ] =      8;
		rom[ 1800 ] =      0;
		rom[ 1801 ] =    -87;
		rom[ 1802 ] =     38;
		rom[ 1803 ] =      7;
		rom[ 1804 ] =     47;
		rom[ 1805 ] =     20;
		rom[ 1806 ] =     57;
		rom[ 1807 ] =     16;
		rom[ 1808 ] =     56;
		rom[ 1809 ] =   -111;
		rom[ 1810 ] =     97;
		rom[ 1811 ] =    102;
		rom[ 1812 ] =    -68;
		rom[ 1813 ] =    -17;
		rom[ 1814 ] =     40;
		rom[ 1815 ] =    198;
		rom[ 1816 ] =   -154;
		rom[ 1817 ] =   -158;
		rom[ 1818 ] =   -181;
		rom[ 1819 ] =    -18;
		rom[ 1820 ] =     21;
		rom[ 1821 ] =     70;
		rom[ 1822 ] =    -15;
		rom[ 1823 ] =    -15;
		rom[ 1824 ] =    129;
		rom[ 1825 ] =     78;
		rom[ 1826 ] =   -128;
		rom[ 1827 ] =    100;
		rom[ 1828 ] =     51;
		rom[ 1829 ] =   -136;
		rom[ 1830 ] =   -160;
		rom[ 1831 ] =    363;
		rom[ 1832 ] =     40;
		rom[ 1833 ] =    -42;
		rom[ 1834 ] =     38;
		rom[ 1835 ] =    108;
		rom[ 1836 ] =     37;
		rom[ 1837 ] =     68;
		rom[ 1838 ] =    110;
		rom[ 1839 ] =    177;
		rom[ 1840 ] =    -86;
		rom[ 1841 ] =   -346;
		rom[ 1842 ] =    -15;
		rom[ 1843 ] =    -10;
		rom[ 1844 ] =     60;
		rom[ 1845 ] =    -54;
		rom[ 1846 ] =     53;
		rom[ 1847 ] =     -2;
		rom[ 1848 ] =     11;
		rom[ 1849 ] =    -60;
		rom[ 1850 ] =     70;
		rom[ 1851 ] =     19;
		rom[ 1852 ] =     -5;
		rom[ 1853 ] =    -10;
		rom[ 1854 ] =    128;
		rom[ 1855 ] =     67;
		rom[ 1856 ] =     81;
		rom[ 1857 ] =    -35;
		rom[ 1858 ] =     -7;
		rom[ 1859 ] =     -3;
		rom[ 1860 ] =     11;
		rom[ 1861 ] =     81;
		rom[ 1862 ] =     43;
		rom[ 1863 ] =    -37;
		rom[ 1864 ] =     31;
		rom[ 1865 ] =     -6;
		rom[ 1866 ] =     42;
		rom[ 1867 ] =    288;
		rom[ 1868 ] =      9;
		rom[ 1869 ] =    -52;
		rom[ 1870 ] =    138;
		rom[ 1871 ] =      0;
		rom[ 1872 ] =    107;
		rom[ 1873 ] =     32;
		rom[ 1874 ] =     55;
		rom[ 1875 ] =   -105;
		rom[ 1876 ] =     28;
		rom[ 1877 ] =    -76;
		rom[ 1878 ] =     63;
		rom[ 1879 ] =    -59;
		rom[ 1880 ] =     39;
		rom[ 1881 ] =    -13;
		rom[ 1882 ] =   -595;
		rom[ 1883 ] =     -2;
		rom[ 1884 ] =   -171;
		rom[ 1885 ] =   -324;
		rom[ 1886 ] =      3;
		rom[ 1887 ] =     -6;
		rom[ 1888 ] =     -7;
		rom[ 1889 ] =    -36;
		rom[ 1890 ] =     96;
		rom[ 1891 ] =   -867;
		rom[ 1892 ] =      4;
		rom[ 1893 ] =    -45;
		rom[ 1894 ] =    -79;
		rom[ 1895 ] =     84;
		rom[ 1896 ] =    -46;
		rom[ 1897 ] =   -289;
		rom[ 1898 ] =     17;
		rom[ 1899 ] =     -4;
		rom[ 1900 ] =    -47;
		rom[ 1901 ] =     -4;
		rom[ 1902 ] =      3;
		rom[ 1903 ] =   -106;
		rom[ 1904 ] =     30;
		rom[ 1905 ] =    -50;
		rom[ 1906 ] =     -6;
		rom[ 1907 ] =     -6;
		rom[ 1908 ] =     16;
		rom[ 1909 ] =      0;
		rom[ 1910 ] =    125;
		rom[ 1911 ] =    130;
		rom[ 1912 ] =    -41;
		rom[ 1913 ] =   -289;
		rom[ 1914 ] =     22;
		rom[ 1915 ] =    -37;
		rom[ 1916 ] =    219;
		rom[ 1917 ] =     86;
		rom[ 1918 ] =     30;
		rom[ 1919 ] =    -62;
		rom[ 1920 ] =    -75;
		rom[ 1921 ] =      0;
		rom[ 1922 ] =    -36;
		rom[ 1923 ] =    -72;
		rom[ 1924 ] =    -72;
		rom[ 1925 ] =    156;
		rom[ 1926 ] =   -105;
		rom[ 1927 ] =     75;
		rom[ 1928 ] =     36;
		rom[ 1929 ] =   -175;
		rom[ 1930 ] =     31;
		rom[ 1931 ] =   -262;
		rom[ 1932 ] =     54;
		rom[ 1933 ] =    124;
		rom[ 1934 ] =     80;
		rom[ 1935 ] =    -76;
		rom[ 1936 ] =   -255;
		rom[ 1937 ] =      5;
		rom[ 1938 ] =     -7;
		rom[ 1939 ] =    -68;
		rom[ 1940 ] =    -96;
		rom[ 1941 ] =    105;
		rom[ 1942 ] =     33;
		rom[ 1943 ] =      0;
		rom[ 1944 ] =    -54;
		rom[ 1945 ] =     -2;
		rom[ 1946 ] =    -14;
		rom[ 1947 ] =   -187;
		rom[ 1948 ] =     42;
		rom[ 1949 ] =   -238;
		rom[ 1950 ] =     64;
		rom[ 1951 ] =     17;
		rom[ 1952 ] =     41;
		rom[ 1953 ] =     -5;
		rom[ 1954 ] =    -39;
		rom[ 1955 ] =    188;
		rom[ 1956 ] =     46;
		rom[ 1957 ] =     -3;
		rom[ 1958 ] =     -9;
		rom[ 1959 ] =    108;
		rom[ 1960 ] =   -252;
		rom[ 1961 ] =     54;
		rom[ 1962 ] =     76;
		rom[ 1963 ] =    -62;
		rom[ 1964 ] =     36;
		rom[ 1965 ] =    -52;
		rom[ 1966 ] =    102;
		rom[ 1967 ] =    -13;
		rom[ 1968 ] =    318;
		rom[ 1969 ] =    153;
		rom[ 1970 ] =     40;
		rom[ 1971 ] =   -116;
		rom[ 1972 ] =     57;
		rom[ 1973 ] =    -61;
		rom[ 1974 ] =     10;
		rom[ 1975 ] =     36;
		rom[ 1976 ] =     21;
		rom[ 1977 ] =     -8;
		rom[ 1978 ] =     13;
		rom[ 1979 ] =    -86;
		rom[ 1980 ] =   -104;
		rom[ 1981 ] =   -209;
		rom[ 1982 ] =    -83;
		rom[ 1983 ] =     11;
		rom[ 1984 ] =     56;
		rom[ 1985 ] =    -56;
		rom[ 1986 ] =     45;
		rom[ 1987 ] =   -223;
		rom[ 1988 ] =      5;
		rom[ 1989 ] =     13;
		rom[ 1990 ] =     88;
		rom[ 1991 ] =   -167;
		rom[ 1992 ] =    150;
		rom[ 1993 ] =    -82;
		rom[ 1994 ] =    -60;
		rom[ 1995 ] =   -411;
		rom[ 1996 ] =     38;
		rom[ 1997 ] =      3;
		rom[ 1998 ] =    142;
		rom[ 1999 ] =    -96;
		rom[ 2000 ] =   -109;
		rom[ 2001 ] =     11;
		rom[ 2002 ] =     11;
		rom[ 2003 ] =    -45;
		rom[ 2004 ] =    -76;
		rom[ 2005 ] =    -12;
		rom[ 2006 ] =     47;
		rom[ 2007 ] =    -46;
		rom[ 2008 ] =    -16;
		rom[ 2009 ] =    -15;
		rom[ 2010 ] =   -361;
		rom[ 2011 ] =    -13;
		rom[ 2012 ] =    113;
		rom[ 2013 ] =    -47;
		rom[ 2014 ] =    208;
		rom[ 2015 ] =      0;
		rom[ 2016 ] =     14;
		rom[ 2017 ] =    -51;
		rom[ 2018 ] =     58;
		rom[ 2019 ] =    -66;
		rom[ 2020 ] =     33;
		rom[ 2021 ] =      4;
		rom[ 2022 ] =     36;
		rom[ 2023 ] =   -143;
		rom[ 2024 ] =    -75;
		rom[ 2025 ] =      3;
		rom[ 2026 ] =      0;
		rom[ 2027 ] =    -10;
		rom[ 2028 ] =    -64;
		rom[ 2029 ] =    -46;
		rom[ 2030 ] =     37;
		rom[ 2031 ] =     87;
		rom[ 2032 ] =   -258;
		rom[ 2033 ] =     21;
		rom[ 2034 ] =     15;
		rom[ 2035 ] =     21;
		rom[ 2036 ] =     30;
		rom[ 2037 ] =    486;
		rom[ 2038 ] =     66;
		rom[ 2039 ] =     11;
		rom[ 2040 ] =    -10;
		rom[ 2041 ] =    -18;
		rom[ 2042 ] =    220;
		rom[ 2043 ] =    -40;
		rom[ 2044 ] =   -654;
		rom[ 2045 ] =   -181;
		rom[ 2046 ] =    422;
		rom[ 2047 ] =    -44;
		rom[ 2048 ] =    -20;
		rom[ 2049 ] =     25;
		rom[ 2050 ] =     68;
		rom[ 2051 ] =   -217;
		rom[ 2052 ] =   -143;
		rom[ 2053 ] =    248;
		rom[ 2054 ] =   -281;
		rom[ 2055 ] =    210;
		rom[ 2056 ] =     73;
		rom[ 2057 ] =   -200;
		rom[ 2058 ] =     52;
		rom[ 2059 ] =     16;
		rom[ 2060 ] =    -45;
		rom[ 2061 ] =    283;
		rom[ 2062 ] =    178;
		rom[ 2063 ] =    -64;
		rom[ 2064 ] =     29;
		rom[ 2065 ] =    -13;
		rom[ 2066 ] =     11;
		rom[ 2067 ] =    -88;
		rom[ 2068 ] =     29;
		rom[ 2069 ] =   -112;
		rom[ 2070 ] =   -186;
		rom[ 2071 ] =    -46;
		rom[ 2072 ] =      9;
		rom[ 2073 ] =    -53;
		rom[ 2074 ] =     71;
		rom[ 2075 ] =    139;
		rom[ 2076 ] =    -28;
		rom[ 2077 ] =    -42;
		rom[ 2078 ] =   -201;
		rom[ 2079 ] =    170;
		rom[ 2080 ] =     41;
		rom[ 2081 ] =    -40;
		rom[ 2082 ] =  -1149;
		rom[ 2083 ] =      3;
		rom[ 2084 ] =     33;
		rom[ 2085 ] =   -187;
		rom[ 2086 ] =     35;
		rom[ 2087 ] =     20;
		rom[ 2088 ] =    107;
		rom[ 2089 ] =    165;
		rom[ 2090 ] =     36;
		rom[ 2091 ] =   -599;
		rom[ 2092 ] =     21;
		rom[ 2093 ] =    -13;
		rom[ 2094 ] =    188;
		rom[ 2095 ] =    178;
		rom[ 2096 ] =    -52;
		rom[ 2097 ] =    -45;
		rom[ 2098 ] =     48;
		rom[ 2099 ] =    839;
		rom[ 2100 ] =     60;
		rom[ 2101 ] =     76;
		rom[ 2102 ] =    -34;
		rom[ 2103 ] =    -74;
		rom[ 2104 ] =   -174;
		rom[ 2105 ] =     -3;
		rom[ 2106 ] =    278;
		rom[ 2107 ] =     50;
		rom[ 2108 ] =   -145;
		rom[ 2109 ] =     36;
		rom[ 2110 ] =   -142;
		rom[ 2111 ] =    -58;
		rom[ 2112 ] =     50;
		rom[ 2113 ] =    -87;
		rom[ 2114 ] =     23;
		rom[ 2115 ] =      0;
		rom[ 2116 ] =      6;
		rom[ 2117 ] =    -12;
		rom[ 2118 ] =   -131;
		rom[ 2119 ] =   -305;
		rom[ 2120 ] =      9;
		rom[ 2121 ] =    126;
		rom[ 2122 ] =    102;
		rom[ 2123 ] =    176;
		rom[ 2124 ] =     65;
		rom[ 2125 ] =     79;
		rom[ 2126 ] =    -70;
		rom[ 2127 ] =    -69;
		rom[ 2128 ] =   -226;
		rom[ 2129 ] =   -139;
		rom[ 2130 ] =      6;
		rom[ 2131 ] =     54;
		rom[ 2132 ] =   -174;
		rom[ 2133 ] =     60;
		rom[ 2134 ] =    -54;
		rom[ 2135 ] =    172;
		rom[ 2136 ] =   -206;
		rom[ 2137 ] =      4;
		rom[ 2138 ] =    120;
		rom[ 2139 ] =    -15;
		rom[ 2140 ] =   -260;
		rom[ 2141 ] =      1;
		rom[ 2142 ] =      0;
		rom[ 2143 ] =     63;
		rom[ 2144 ] =   -240;
		rom[ 2145 ] =      2;
		rom[ 2146 ] =    -91;
		rom[ 2147 ] =   -417;
		rom[ 2148 ] =   -434;
		rom[ 2149 ] =    132;
		rom[ 2150 ] =    243;
		rom[ 2151 ] =   -296;
		rom[ 2152 ] =    -84;
		rom[ 2153 ] =      0;
		rom[ 2154 ] =   -198;
		rom[ 2155 ] =    190;
		rom[ 2156 ] =    -47;
		rom[ 2157 ] =      8;
		rom[ 2158 ] =   -327;
		rom[ 2159 ] =    170;
		rom[ 2160 ] =     -5;
		rom[ 2161 ] =     59;
		rom[ 2162 ] =    219;
		rom[ 2163 ] =      7;
		rom[ 2164 ] =   -247;
		rom[ 2165 ] =    132;
		rom[ 2166 ] =    -46;
		rom[ 2167 ] =     81;
		rom[ 2168 ] =    -15;
		rom[ 2169 ] =      5;
		rom[ 2170 ] =    -74;
		rom[ 2171 ] =     59;
		rom[ 2172 ] =    -66;
		rom[ 2173 ] =     15;
		rom[ 2174 ] =    419;
		rom[ 2175 ] =   -114;
		rom[ 2176 ] =    -60;
		rom[ 2177 ] =    206;
		rom[ 2178 ] =    -84;
		rom[ 2179 ] =   -363;
		rom[ 2180 ] =    149;
		rom[ 2181 ] =     99;
		rom[ 2182 ] =    -40;
		rom[ 2183 ] =      2;
		rom[ 2184 ] =     -8;
		rom[ 2185 ] =     41;
		rom[ 2186 ] =    139;
		rom[ 2187 ] =     -3;
		rom[ 2188 ] =    194;
		rom[ 2189 ] =   -189;
		rom[ 2190 ] =    393;
		rom[ 2191 ] =     52;
		rom[ 2192 ] =     13;
		rom[ 2193 ] =     75;
		rom[ 2194 ] =    -72;
		rom[ 2195 ] =     22;
		rom[ 2196 ] =     64;
		rom[ 2197 ] =      4;
		rom[ 2198 ] =    -64;
		rom[ 2199 ] =     22;
		rom[ 2200 ] =   -104;
		rom[ 2201 ] =     44;
		rom[ 2202 ] =     -9;
		rom[ 2203 ] =   -206;
		rom[ 2204 ] =    -44;
		rom[ 2205 ] =   -503;
		rom[ 2206 ] =   -263;
		rom[ 2207 ] =     31;
		rom[ 2208 ] =    190;
		rom[ 2209 ] =   -113;
		rom[ 2210 ] =    -44;
		rom[ 2211 ] =    -31;
		rom[ 2212 ] =    -85;
		rom[ 2213 ] =     37;
		rom[ 2214 ] =     -7;
		rom[ 2215 ] =     84;
		rom[ 2216 ] =   -213;
		rom[ 2217 ] =     45;
		rom[ 2218 ] =     17;
		rom[ 2219 ] =    -96;
		rom[ 2220 ] =    -53;
		rom[ 2221 ] =    116;
		rom[ 2222 ] =     19;
		rom[ 2223 ] =    -72;
		rom[ 2224 ] =   -141;
		rom[ 2225 ] =    -53;
		rom[ 2226 ] =     17;
		rom[ 2227 ] =    193;
		rom[ 2228 ] =    -81;
		rom[ 2229 ] =   -291;
		rom[ 2230 ] =     48;
		rom[ 2231 ] =     42;
		rom[ 2232 ] =     -5;
		rom[ 2233 ] =    135;
		rom[ 2234 ] =    -71;
		rom[ 2235 ] =     16;
		rom[ 2236 ] =    130;
		rom[ 2237 ] =   -371;
		rom[ 2238 ] =      6;
		rom[ 2239 ] =     30;
		rom[ 2240 ] =   -261;
		rom[ 2241 ] =     47;
		rom[ 2242 ] =   -212;
		rom[ 2243 ] =     36;
		rom[ 2244 ] =    122;
		rom[ 2245 ] =   -156;
		rom[ 2246 ] =     30;
		rom[ 2247 ] =     16;
		rom[ 2248 ] =    -36;
		rom[ 2249 ] =     16;
		rom[ 2250 ] =   -138;
		rom[ 2251 ] =    100;
		rom[ 2252 ] =   -138;
		rom[ 2253 ] =      9;
		rom[ 2254 ] =    586;
		rom[ 2255 ] =   -153;
		rom[ 2256 ] =     95;
		rom[ 2257 ] =     12;
		rom[ 2258 ] =    -18;
		rom[ 2259 ] =    -11;
		rom[ 2260 ] =   -204;
		rom[ 2261 ] =   -161;
		rom[ 2262 ] =    -10;
		rom[ 2263 ] =   -404;
		rom[ 2264 ] =    -12;
		rom[ 2265 ] =     -8;
		rom[ 2266 ] =     43;
		rom[ 2267 ] =     41;
		rom[ 2268 ] =    144;
		rom[ 2269 ] =     30;
		rom[ 2270 ] =    237;
		rom[ 2271 ] =    -41;
		rom[ 2272 ] =    260;
		rom[ 2273 ] =      8;
		rom[ 2274 ] =     -2;
		rom[ 2275 ] =    -29;
		rom[ 2276 ] =    -17;
		rom[ 2277 ] =   -172;
		rom[ 2278 ] =   -190;
		rom[ 2279 ] =     -6;
		rom[ 2280 ] =    -54;
		rom[ 2281 ] =     36;
		rom[ 2282 ] =    -17;
		rom[ 2283 ] =   -579;
		rom[ 2284 ] =    -38;
		rom[ 2285 ] =    106;
		rom[ 2286 ] =   -106;
		rom[ 2287 ] =     15;
		rom[ 2288 ] =    118;
		rom[ 2289 ] =   -338;
		rom[ 2290 ] =     49;
		rom[ 2291 ] =     19;
		rom[ 2292 ] =    117;
		rom[ 2293 ] =   -127;
		rom[ 2294 ] =   -394;
		rom[ 2295 ] =     29;
		rom[ 2296 ] =   -375;
		rom[ 2297 ] =    -28;
		rom[ 2298 ] =    146;
		rom[ 2299 ] =     24;
		rom[ 2300 ] =    222;
		rom[ 2301 ] =     14;
		rom[ 2302 ] =    -71;
		rom[ 2303 ] =     75;
		rom[ 2304 ] =    155;
		rom[ 2305 ] =    100;
		rom[ 2306 ] =    150;
		rom[ 2307 ] =    163;
		rom[ 2308 ] =    -37;
		rom[ 2309 ] =    -74;
		rom[ 2310 ] =    134;
		rom[ 2311 ] =   -228;
		rom[ 2312 ] =    113;
		rom[ 2313 ] =     45;
		rom[ 2314 ] =    -76;
		rom[ 2315 ] =    409;
		rom[ 2316 ] =   -136;
		rom[ 2317 ] =   -107;
		rom[ 2318 ] =     33;
		rom[ 2319 ] =    251;
		rom[ 2320 ] =   -144;
		rom[ 2321 ] =     -2;
		rom[ 2322 ] =     34;
		rom[ 2323 ] =     24;
		rom[ 2324 ] =    -10;
		rom[ 2325 ] =     -7;
		rom[ 2326 ] =     57;
		rom[ 2327 ] =     -7;
		rom[ 2328 ] =     32;
		rom[ 2329 ] =     65;
		rom[ 2330 ] =     39;
		rom[ 2331 ] =      0;
		rom[ 2332 ] =   -141;
		rom[ 2333 ] =    -44;
		rom[ 2334 ] =     10;
		rom[ 2335 ] =     -3;
		rom[ 2336 ] =     -4;
		rom[ 2337 ] =     35;
		rom[ 2338 ] =     60;
		rom[ 2339 ] =   -331;
		rom[ 2340 ] =    -47;
		rom[ 2341 ] =    -50;
		rom[ 2342 ] =    -83;
		rom[ 2343 ] =     -1;
		rom[ 2344 ] =    151;
		rom[ 2345 ] =    -60;
		rom[ 2346 ] =    187;
		rom[ 2347 ] =    279;
		rom[ 2348 ] =     43;
		rom[ 2349 ] =    257;
		rom[ 2350 ] =    -13;
		rom[ 2351 ] =   -240;
		rom[ 2352 ] =    139;
		rom[ 2353 ] =    103;
		rom[ 2354 ] =      8;
		rom[ 2355 ] =    -89;
		rom[ 2356 ] =     43;
		rom[ 2357 ] =    -51;
		rom[ 2358 ] =   -126;
		rom[ 2359 ] =     -4;
		rom[ 2360 ] =    -42;
		rom[ 2361 ] =   -106;
		rom[ 2362 ] =    181;
		rom[ 2363 ] =    -78;
		rom[ 2364 ] =      6;
		rom[ 2365 ] =    -42;
		rom[ 2366 ] =     51;
		rom[ 2367 ] =      1;
		rom[ 2368 ] =    224;
		rom[ 2369 ] =    -44;
		rom[ 2370 ] =   -155;
		rom[ 2371 ] =    -49;
		rom[ 2372 ] =     41;
		rom[ 2373 ] =   -196;
		rom[ 2374 ] =    -29;
		rom[ 2375 ] =     -9;
		rom[ 2376 ] =     47;
		rom[ 2377 ] =      1;
		rom[ 2378 ] =     31;
		rom[ 2379 ] =    -49;
		rom[ 2380 ] =     62;
		rom[ 2381 ] =    -99;
		rom[ 2382 ] =  -7680;
		rom[ 2383 ] =    -16;
		rom[ 2384 ] =   -179;
		rom[ 2385 ] =     15;
		rom[ 2386 ] =      0;
		rom[ 2387 ] =    -36;
		rom[ 2388 ] =      0;
		rom[ 2389 ] =     -4;
		rom[ 2390 ] =   -107;
		rom[ 2391 ] =    -52;
		rom[ 2392 ] =     45;
		rom[ 2393 ] =      7;
		rom[ 2394 ] =     77;
		rom[ 2395 ] =    -67;
		rom[ 2396 ] =     18;
		rom[ 2397 ] =   -219;
		rom[ 2398 ] =    -12;
		rom[ 2399 ] =   -115;
		rom[ 2400 ] =   -119;
		rom[ 2401 ] =    -11;
		rom[ 2402 ] =     73;
		rom[ 2403 ] =     -2;
		rom[ 2404 ] =   -902;
		rom[ 2405 ] =    375;
		rom[ 2406 ] =   -333;
		rom[ 2407 ] =     -2;
		rom[ 2408 ] =     21;
		rom[ 2409 ] =    -43;
		rom[ 2410 ] =     64;
		rom[ 2411 ] =    -62;
		rom[ 2412 ] =     51;
		rom[ 2413 ] =   -272;
		rom[ 2414 ] =    127;
		rom[ 2415 ] =    106;
		rom[ 2416 ] =     34;
		rom[ 2417 ] =    149;
		rom[ 2418 ] =   -805;
		rom[ 2419 ] =    177;
		rom[ 2420 ] =     77;
		rom[ 2421 ] =    -81;
		rom[ 2422 ] =     14;
		rom[ 2423 ] =    235;
		rom[ 2424 ] =     51;
		rom[ 2425 ] =      5;
		rom[ 2426 ] =     33;
		rom[ 2427 ] =    -49;
		rom[ 2428 ] =     40;
		rom[ 2429 ] =   -141;
		rom[ 2430 ] =    -11;
		rom[ 2431 ] =   -241;
		rom[ 2432 ] =     -1;
		rom[ 2433 ] =     -5;
		rom[ 2434 ] =     28;
		rom[ 2435 ] =      2;
		rom[ 2436 ] =    -21;
		rom[ 2437 ] =    290;
		rom[ 2438 ] =    195;
		rom[ 2439 ] =    -15;
		rom[ 2440 ] =     23;
		rom[ 2441 ] =     21;
		rom[ 2442 ] =   -281;
		rom[ 2443 ] =    -51;
		rom[ 2444 ] =     36;
		rom[ 2445 ] =   -315;
		rom[ 2446 ] =      3;
		rom[ 2447 ] =    -82;
		rom[ 2448 ] =     58;
		rom[ 2449 ] =    130;
		rom[ 2450 ] =     18;
		rom[ 2451 ] =     40;
		rom[ 2452 ] =    -45;
		rom[ 2453 ] =     14;
		rom[ 2454 ] =    -18;
		rom[ 2455 ] =    -50;
		rom[ 2456 ] =   -220;
		rom[ 2457 ] =   -290;
		rom[ 2458 ] =     40;
		rom[ 2459 ] =   -157;
		rom[ 2460 ] =    178;
		rom[ 2461 ] =    -38;
		rom[ 2462 ] =     44;
		rom[ 2463 ] =    158;
		rom[ 2464 ] =    108;
		rom[ 2465 ] =    320;
		rom[ 2466 ] =     36;
		rom[ 2467 ] =    152;
		rom[ 2468 ] =   -201;
		rom[ 2469 ] =   -364;
		rom[ 2470 ] =      7;
		rom[ 2471 ] =    -57;
		rom[ 2472 ] =     81;
		rom[ 2473 ] =    166;
		rom[ 2474 ] =     28;
		rom[ 2475 ] =      5;
		rom[ 2476 ] =      8;
		rom[ 2477 ] =    -65;
		rom[ 2478 ] =    232;
		rom[ 2479 ] =      2;
		rom[ 2480 ] =   -245;
		rom[ 2481 ] =    350;
		rom[ 2482 ] =     55;
		rom[ 2483 ] =   -226;
		rom[ 2484 ] =     16;
		rom[ 2485 ] =    -38;
		rom[ 2486 ] =     32;
		rom[ 2487 ] =    -16;
		rom[ 2488 ] =     28;
		rom[ 2489 ] =     93;
		rom[ 2490 ] =     70;
		rom[ 2491 ] =    276;
		rom[ 2492 ] =     52;
		rom[ 2493 ] =      6;
		rom[ 2494 ] =     14;
		rom[ 2495 ] =     53;
		rom[ 2496 ] =   -400;
		rom[ 2497 ] =    134;
		rom[ 2498 ] =   -335;
		rom[ 2499 ] =   -130;
		rom[ 2500 ] =     16;
		rom[ 2501 ] =    787;
		rom[ 2502 ] =     99;
		rom[ 2503 ] =    115;
		rom[ 2504 ] =    109;
		rom[ 2505 ] =   -170;
		rom[ 2506 ] =     71;
		rom[ 2507 ] =    113;
		rom[ 2508 ] =    -64;
		rom[ 2509 ] =     88;
		rom[ 2510 ] =      8;
		rom[ 2511 ] =    -15;
		rom[ 2512 ] =    -62;
		rom[ 2513 ] =   -123;
		rom[ 2514 ] =    184;
		rom[ 2515 ] =    -87;
		rom[ 2516 ] =   -210;
		rom[ 2517 ] =     48;
		rom[ 2518 ] =     -7;
		rom[ 2519 ] =   -138;
		rom[ 2520 ] =    -10;
		rom[ 2521 ] =     39;
		rom[ 2522 ] =    -56;
		rom[ 2523 ] =    155;
		rom[ 2524 ] =     -3;
		rom[ 2525 ] =    -70;
		rom[ 2526 ] =    -10;
		rom[ 2527 ] =    -14;
		rom[ 2528 ] =   -140;
		rom[ 2529 ] =    123;
		rom[ 2530 ] =    -84;
		rom[ 2531 ] =     32;
		rom[ 2532 ] =    138;
		rom[ 2533 ] =     11;
		rom[ 2534 ] =    106;
		rom[ 2535 ] =    176;
		rom[ 2536 ] =    -58;
		rom[ 2537 ] =    -55;
		rom[ 2538 ] =   -185;
		rom[ 2539 ] =     47;
		rom[ 2540 ] =   -118;
		rom[ 2541 ] =     61;
		rom[ 2542 ] =      8;
		rom[ 2543 ] =     19;
		rom[ 2544 ] =    -47;
		rom[ 2545 ] =  -7680;
		rom[ 2546 ] =    -12;
		rom[ 2547 ] =     40;
		rom[ 2548 ] =    -64;
		rom[ 2549 ] =     47;
		rom[ 2550 ] =    -49;
		rom[ 2551 ] =     58;
		rom[ 2552 ] =   -170;
		rom[ 2553 ] =    165;
		rom[ 2554 ] =     89;
		rom[ 2555 ] =     53;
		rom[ 2556 ] =    -45;
		rom[ 2557 ] =     78;
		rom[ 2558 ] =    256;
		rom[ 2559 ] =    -16;
		rom[ 2560 ] =    -78;
		rom[ 2561 ] =   -240;
		rom[ 2562 ] =     -6;
		rom[ 2563 ] =     21;
		rom[ 2564 ] =    -79;
		rom[ 2565 ] =   -216;
		rom[ 2566 ] =   -342;
		rom[ 2567 ] =   -155;
		rom[ 2568 ] =     -9;
		rom[ 2569 ] =     83;
		rom[ 2570 ] =     75;
		rom[ 2571 ] =   -384;
		rom[ 2572 ] =    -11;
		rom[ 2573 ] =    -37;
		rom[ 2574 ] =     -9;
		rom[ 2575 ] =    153;
		rom[ 2576 ] =     -9;
		rom[ 2577 ] =     14;
		rom[ 2578 ] =    -67;
		rom[ 2579 ] =     91;
		rom[ 2580 ] =    131;
		rom[ 2581 ] =      0;
		rom[ 2582 ] =    157;
		rom[ 2583 ] =     46;
		rom[ 2584 ] =   -493;
		rom[ 2585 ] =    157;
		rom[ 2586 ] =    113;
		rom[ 2587 ] =     62;
		rom[ 2588 ] =    -38;
		rom[ 2589 ] =    -46;
		rom[ 2590 ] =    -48;
		rom[ 2591 ] =     58;
		rom[ 2592 ] =   -132;
		rom[ 2593 ] =     89;
		rom[ 2594 ] =    -55;
		rom[ 2595 ] =    -73;
		rom[ 2596 ] =     67;
		rom[ 2597 ] =   -127;
		rom[ 2598 ] =   -197;
		rom[ 2599 ] =    -82;
		rom[ 2600 ] =    -57;
		rom[ 2601 ] =    131;
		rom[ 2602 ] =     12;
		rom[ 2603 ] =      1;
		rom[ 2604 ] =     17;
		rom[ 2605 ] =   -485;
		rom[ 2606 ] =   -365;
		rom[ 2607 ] =     46;
		rom[ 2608 ] =    -42;
		rom[ 2609 ] =    -71;
		rom[ 2610 ] =     -4;
		rom[ 2611 ] =     -1;
		rom[ 2612 ] =    650;
		rom[ 2613 ] =     73;
		rom[ 2614 ] =    167;
		rom[ 2615 ] =     69;
		rom[ 2616 ] =    -64;
		rom[ 2617 ] =     14;
		rom[ 2618 ] =    119;
		rom[ 2619 ] =     65;
		rom[ 2620 ] =     18;
		rom[ 2621 ] =     43;
		rom[ 2622 ] =    -45;
		rom[ 2623 ] =    611;
		rom[ 2624 ] =    159;
		rom[ 2625 ] =    -16;
		rom[ 2626 ] =     27;
		rom[ 2627 ] =   -234;
		rom[ 2628 ] =    381;
		rom[ 2629 ] =     50;
		rom[ 2630 ] =      0;
		rom[ 2631 ] =    267;
		rom[ 2632 ] =     69;
		rom[ 2633 ] =     14;
		rom[ 2634 ] =   -247;
		rom[ 2635 ] =    -89;
		rom[ 2636 ] =    -13;
		rom[ 2637 ] =     71;
		rom[ 2638 ] =     53;
		rom[ 2639 ] =     29;
		rom[ 2640 ] =    -57;
		rom[ 2641 ] =    -25;
		rom[ 2642 ] =     20;
		rom[ 2643 ] =     41;
		rom[ 2644 ] =    -44;
		rom[ 2645 ] =     32;
		rom[ 2646 ] =   -284;
		rom[ 2647 ] =  -1234;
		rom[ 2648 ] =   -163;
		rom[ 2649 ] =    628;
		rom[ 2650 ] =   -130;
		rom[ 2651 ] =     28;
		rom[ 2652 ] =   -362;
		rom[ 2653 ] =     10;
		rom[ 2654 ] =     85;
		rom[ 2655 ] =     11;
		rom[ 2656 ] =      0;
		rom[ 2657 ] =     91;
		rom[ 2658 ] =    112;
		rom[ 2659 ] =    -11;
		rom[ 2660 ] =   -235;
		rom[ 2661 ] =     51;
		rom[ 2662 ] =    -59;
		rom[ 2663 ] =     68;
		rom[ 2664 ] =     12;
		rom[ 2665 ] =   -724;
		rom[ 2666 ] =    -40;
		rom[ 2667 ] =   -510;
		rom[ 2668 ] =    334;
		rom[ 2669 ] =    -11;
		rom[ 2670 ] =    -52;
		rom[ 2671 ] =   -244;
		rom[ 2672 ] =   -541;
		rom[ 2673 ] =   -412;
		rom[ 2674 ] =    179;
		rom[ 2675 ] =   -102;
		rom[ 2676 ] =    113;
		rom[ 2677 ] =   -403;
		rom[ 2678 ] =    -10;
		rom[ 2679 ] =     -3;
		rom[ 2680 ] =      6;
		rom[ 2681 ] =    -16;
		rom[ 2682 ] =   -215;
		rom[ 2683 ] =     41;
		rom[ 2684 ] =      1;
		rom[ 2685 ] =     34;
		rom[ 2686 ] =    -41;
		rom[ 2687 ] =    141;
		rom[ 2688 ] =   -275;
		rom[ 2689 ] =    299;
		rom[ 2690 ] =     97;
		rom[ 2691 ] =     28;
		rom[ 2692 ] =    -47;
		rom[ 2693 ] =     47;
		rom[ 2694 ] =    243;
		rom[ 2695 ] =      9;
		rom[ 2696 ] =    -16;
		rom[ 2697 ] =    107;
		rom[ 2698 ] =    -54;
		rom[ 2699 ] =   -544;
		rom[ 2700 ] =   -380;
		rom[ 2701 ] =     82;
		rom[ 2702 ] =     48;
		rom[ 2703 ] =     71;
		rom[ 2704 ] =     68;
		rom[ 2705 ] =   -155;
		rom[ 2706 ] =      5;
		rom[ 2707 ] =    124;
		rom[ 2708 ] =   -238;
		rom[ 2709 ] =     87;
		rom[ 2710 ] =    -15;
		rom[ 2711 ] =    164;
		rom[ 2712 ] =   -101;
		rom[ 2713 ] =   -117;
		rom[ 2714 ] =     55;
		rom[ 2715 ] =    108;
		rom[ 2716 ] =   -162;
		rom[ 2717 ] =    -77;
		rom[ 2718 ] =    103;
		rom[ 2719 ] =   -199;
		rom[ 2720 ] =     41;
		rom[ 2721 ] =   -204;
		rom[ 2722 ] =     65;
		rom[ 2723 ] =   -181;
		rom[ 2724 ] =    189;
		rom[ 2725 ] =    -62;
		rom[ 2726 ] =    -33;
		rom[ 2727 ] =     35;
		rom[ 2728 ] =    229;
		rom[ 2729 ] =   -220;
		rom[ 2730 ] =    218;
		rom[ 2731 ] =    -75;
		rom[ 2732 ] =     49;
		rom[ 2733 ] =    -65;
		rom[ 2734 ] =     55;
		rom[ 2735 ] =    -11;
		rom[ 2736 ] =     48;
		rom[ 2737 ] =     80;
		rom[ 2738 ] =     42;
		rom[ 2739 ] =   -159;
		rom[ 2740 ] =     49;
		rom[ 2741 ] =     -3;
		rom[ 2742 ] =     -8;
		rom[ 2743 ] =     53;
		rom[ 2744 ] =     47;
		rom[ 2745 ] =     13;
		rom[ 2746 ] =     49;
		rom[ 2747 ] =    244;
		rom[ 2748 ] =     63;
		rom[ 2749 ] =   -419;
		rom[ 2750 ] =    -23;
		rom[ 2751 ] =    -91;
		rom[ 2752 ] =     51;
		rom[ 2753 ] =    -48;
		rom[ 2754 ] =    209;
		rom[ 2755 ] =   -117;
		rom[ 2756 ] =     36;
		rom[ 2757 ] =    -52;
		rom[ 2758 ] =     13;
		rom[ 2759 ] =    -56;
		rom[ 2760 ] =     36;
		rom[ 2761 ] =    458;
		rom[ 2762 ] =   -483;
		rom[ 2763 ] =    -14;
		rom[ 2764 ] =    -26;
		rom[ 2765 ] =    -12;
		rom[ 2766 ] =    -23;
		rom[ 2767 ] =   -365;
		rom[ 2768 ] =     82;
		rom[ 2769 ] =     -8;
		rom[ 2770 ] =     -4;
		rom[ 2771 ] =    279;
		rom[ 2772 ] =     79;
		rom[ 2773 ] =   -176;
		rom[ 2774 ] =     -1;
		rom[ 2775 ] =     32;
		rom[ 2776 ] =    100;
		rom[ 2777 ] =    -51;
		rom[ 2778 ] =    232;
		rom[ 2779 ] =    -50;
		rom[ 2780 ] =   -132;
		rom[ 2781 ] =     -8;
		rom[ 2782 ] =     32;
		rom[ 2783 ] =   -162;
		rom[ 2784 ] =     16;
		rom[ 2785 ] =     79;
		rom[ 2786 ] =     43;
		rom[ 2787 ] =     90;
		rom[ 2788 ] =   -190;
		rom[ 2789 ] =    106;
		rom[ 2790 ] =      0;
		rom[ 2791 ] =    -42;
		rom[ 2792 ] =   -133;
		rom[ 2793 ] =      0;
		rom[ 2794 ] =     15;
		rom[ 2795 ] =     37;
		rom[ 2796 ] =     33;
		rom[ 2797 ] =   -350;
		rom[ 2798 ] =     -1;
		rom[ 2799 ] =    -79;
		rom[ 2800 ] =     21;
		rom[ 2801 ] =    -45;
		rom[ 2802 ] =     36;
		rom[ 2803 ] =    -60;
		rom[ 2804 ] =     -5;
		rom[ 2805 ] =     -5;
		rom[ 2806 ] =    118;
		rom[ 2807 ] =    102;
		rom[ 2808 ] =      7;
		rom[ 2809 ] =    111;
		rom[ 2810 ] =     17;
		rom[ 2811 ] =    -53;
		rom[ 2812 ] =     92;
		rom[ 2813 ] =    -39;
		rom[ 2814 ] =     71;
		rom[ 2815 ] =    -93;
		rom[ 2816 ] =    106;
		rom[ 2817 ] =    -43;
		rom[ 2818 ] =   -167;
		rom[ 2819 ] =   -117;
		rom[ 2820 ] =     18;
		rom[ 2821 ] =   -257;
		rom[ 2822 ] =    108;
		rom[ 2823 ] =     67;
		rom[ 2824 ] =   -266;
		rom[ 2825 ] =     -5;
		rom[ 2826 ] =    400;
		rom[ 2827 ] =     37;
		rom[ 2828 ] =      0;
		rom[ 2829 ] =     -9;
		rom[ 2830 ] =   -223;
		rom[ 2831 ] =    152;
		rom[ 2832 ] =    -14;
		rom[ 2833 ] =   -348;
		rom[ 2834 ] =     65;
		rom[ 2835 ] =    -36;
		rom[ 2836 ] =     43;
		rom[ 2837 ] =     73;
		rom[ 2838 ] =     52;
		rom[ 2839 ] =    -39;
		rom[ 2840 ] =     19;
		rom[ 2841 ] =     20;
		rom[ 2842 ] =    -94;
		rom[ 2843 ] =   -236;
		rom[ 2844 ] =     20;
		rom[ 2845 ] =    183;
		rom[ 2846 ] =   -224;
		rom[ 2847 ] =   -151;
		rom[ 2848 ] =    123;
		rom[ 2849 ] =     86;
		rom[ 2850 ] =     80;
		rom[ 2851 ] =     45;
		rom[ 2852 ] =    -75;
		rom[ 2853 ] =    -36;
		rom[ 2854 ] =    142;
		rom[ 2855 ] =    -16;
		rom[ 2856 ] =     50;
		rom[ 2857 ] =     75;
		rom[ 2858 ] =    171;
		rom[ 2859 ] =      0;
		rom[ 2860 ] =     30;
		rom[ 2861 ] =   -129;
		rom[ 2862 ] =    -55;
		rom[ 2863 ] =    -38;
		rom[ 2864 ] =    102;
		rom[ 2865 ] =     29;
		rom[ 2866 ] =     21;
		rom[ 2867 ] =    -48;
		rom[ 2868 ] =     40;
		rom[ 2869 ] =   -273;
		rom[ 2870 ] =     13;
		rom[ 2871 ] =    -15;
		rom[ 2872 ] =    169;
		rom[ 2873 ] =     15;
		rom[ 2874 ] =    -63;
		rom[ 2875 ] =    101;
		rom[ 2876 ] =    -24;
		rom[ 2877 ] =   -117;
		rom[ 2878 ] =     37;
		rom[ 2879 ] =    404;
		rom[ 2880 ] =     19;
		rom[ 2881 ] =    120;
		rom[ 2882 ] =     30;
		rom[ 2883 ] =   -214;
		rom[ 2884 ] =     20;
		rom[ 2885 ] =    -45;
		rom[ 2886 ] =     32;
		rom[ 2887 ] =     69;
		rom[ 2888 ] =   -110;
		rom[ 2889 ] =    150;
		rom[ 2890 ] =     -9;
		rom[ 2891 ] =     -5;
		rom[ 2892 ] =     36;
		rom[ 2893 ] =   -106;
		rom[ 2894 ] =     53;
		rom[ 2895 ] =    162;
		rom[ 2896 ] =   -131;
		rom[ 2897 ] =    -45;
		rom[ 2898 ] =    175;
		rom[ 2899 ] =    -40;
		rom[ 2900 ] =    -62;
		rom[ 2901 ] =   -225;
		rom[ 2902 ] =     45;
		rom[ 2903 ] =    -42;
		rom[ 2904 ] =     88;
		rom[ 2905 ] =    221;
		rom[ 2906 ] =     30;
		rom[ 2907 ] =   -230;
		rom[ 2908 ] =   -277;
		rom[ 2909 ] =     -8;
		rom[ 2910 ] =     55;
		rom[ 2911 ] =    430;
		rom[ 2912 ] =      0;	
	end
endmodule

module strong_thresh_rom(
	input 				clk,
	input		[4:0]	addr,
	output	reg	[11:0]	q
	);
	
	reg					[11:0]	rom [31:0];
	always @(posedge clk) q <= rom[addr];
	initial begin
		rom[   0] = -1290 *0.4  ;
		rom[   1] = -1275 *0.4  ;
		rom[   2] = -1191 *0.4  ;
		rom[   3] = -1140 *0.4  ;
		rom[   4] = -1122 *0.4  ;
		rom[   5] = -1057 *0.4  ;
		rom[   6] = -1029 *0.4  ;
		rom[   7] = -994  *0.4  ;
		rom[   8] = -983  *0.4  ;
		rom[   9] = -933  *0.4  ;
		rom[  10] = -990  *0.4  ;	
		rom[  11] = -951  *0.4  ;	
		rom[  12] = -912  *0.4  ;	
		rom[  13] = -947  *0.4  ;	
		rom[  14] = -877  *0.4  ;	
		rom[  15] = -899  *0.4  ;	
		rom[  16] = -920  *0.4  ;	
		rom[  17] = -868  *0.4  ;	
		rom[  18] = -829  *0.4  ;	
		rom[  19] = -821  *0.4  ;	
		rom[  20] = -839  *0.4  ;	
		rom[  21] = -849  *0.4  ;	
		rom[  22] = -833  *0.4  ;	
		rom[  23] = -862  *0.4  ;	
		rom[  24] = -766  *0.4  ;	
	end

endmodule


module weak_stages_rom(
	input 				clk,
	input		[4:0]	addr,
	output reg	[7:0]	q
	);
	
	reg					[7:0]	rom [31:0];
	always @(posedge clk) q <= rom[addr];
	initial begin
		rom[   0] = 8'd9 ;
		rom[   1] = 8'd16 ;
		rom[   2] = 8'd27 ;
		rom[   3] = 8'd32 ;
		rom[   4] = 8'd52 ;
		rom[   5] = 8'd53 ;
		rom[   6] = 8'd62 ;
		rom[   7] = 8'd72 ;
		rom[   8] = 8'd83 ;
		rom[   9] = 8'd91 ;
		rom[  10] = 8'd99 ;
		rom[  11] = 8'd115;
		rom[  12] = 8'd127;
		rom[  13] = 8'd135;
		rom[  14] = 8'd136;
		rom[  15] = 8'd137;
		rom[  16] = 8'd159;
		rom[  17] = 8'd155;
		rom[  18] = 8'd169;
		rom[  19] = 8'd196;
		rom[  20] = 8'd197;
		rom[  21] = 8'd181;
		rom[  22] = 8'd199;
		rom[  23] = 8'd211;
		rom[  24] = 8'd200;
		rom[  25] = 8'd0;
		rom[  26] = 8'd0;
		rom[  27] = 8'd0;
		rom[  28] = 8'd0;
		rom[  29] = 8'd0;
		rom[  30] = 8'd0;
		rom[  31] = 8'd0;
	end
endmodule


module weak_stages_acc_rom(
	input 				clk,
	input		[4:0]	addr,
	output reg	[11:0]	q
	);
	
	reg					[11:0]	rom [31:0];
	always @(posedge clk) q <= rom[addr];
	initial begin
		rom[   0] = 9	;	
		rom[   1] = 25  ;
		rom[   2] = 52  ;
		rom[   3] = 84  ;
		rom[   4] = 136 ;
		rom[   5] = 189 ;
		rom[   6] = 251 ;
		rom[   7] = 323 ;
		rom[   8] = 406 ;
		rom[   9] = 497 ;
		rom[  10] = 596 ;
		rom[  11] = 711 ;
		rom[  12] = 838 ;
		rom[  13] = 973 ;
		rom[  14] = 1109;
		rom[  15] = 1246;
		rom[  16] = 1405;
		rom[  17] = 1560;
		rom[  18] = 1729;
		rom[  19] = 1925;
		rom[  20] = 2122;
		rom[  21] = 2303;
		rom[  22] = 2502;
		rom[  23] = 2713;
		rom[  24] = 2913;
		rom[  25] = 2913;
		rom[  26] = 2913;
		rom[  27] = 2913;
		rom[  28] = 2913;
		rom[  29] = 2913;
		rom[  30] = 2913;
		rom[  31] = 2913;
	end
endmodule